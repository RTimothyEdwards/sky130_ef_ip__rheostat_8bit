magic
tech sky130A
magscale 1 2
timestamp 1716082924
<< poly >>
rect -414 1402 -272 1431
rect -414 990 -368 1402
rect -318 990 -272 1402
rect -414 974 -272 990
rect -414 366 -272 382
rect -414 -46 -368 366
rect -318 -46 -272 366
rect -414 -76 -272 -46
<< polycont >>
rect -368 990 -318 1402
rect -368 -46 -318 366
<< npolyres >>
rect -414 382 -272 974
<< locali >>
rect -414 1402 -272 1431
rect -414 990 -412 1402
rect -318 990 -272 1402
rect -414 974 -272 990
rect -414 366 -272 382
rect -414 -46 -412 366
rect -318 -46 -272 366
rect -414 -76 -272 -46
<< viali >>
rect -412 990 -368 1402
rect -412 -46 -368 366
<< metal1 >>
rect -425 1402 -354 1431
rect -425 990 -412 1402
rect -368 990 -354 1402
rect -425 974 -354 990
rect -425 366 -354 382
rect -425 -46 -412 366
rect -368 -46 -354 366
rect -425 -76 -354 -46
<< end >>
