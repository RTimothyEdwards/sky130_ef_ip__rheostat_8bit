magic
tech sky130A
magscale 1 2
timestamp 1716082924
<< metal1 >>
rect 261 15219 771 15272
rect 261 15178 328 15219
rect 28 15115 328 15178
rect 704 15170 771 15219
rect 704 15115 876 15170
rect 28 15111 98 15115
rect 36 13244 88 13250
rect 36 13186 88 13192
rect 937 13243 989 13249
rect 937 13185 989 13191
rect -18 1607 38 1724
rect 988 1608 1047 1725
rect -18 45 38 100
rect 938 45 1047 100
<< via1 >>
rect 36 13192 88 13244
rect 937 13191 989 13243
<< metal2 >>
rect 142 13278 717 13330
rect 142 13244 194 13278
rect 30 13192 36 13244
rect 88 13192 194 13244
rect 665 13243 717 13278
rect 665 13191 937 13243
rect 989 13191 995 13243
use dac_3v_cell_dummy  dac_3v_cell_dummy_0
array 0 0 1067 0 9 1507
timestamp 1716082924
transform 1 0 -117 0 1 268
box 99 -275 1166 1410
<< end >>
