VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_ef_ip__rheostat_8bit
  CLASS BLOCK ;
  FOREIGN sky130_ef_ip__rheostat_8bit ;
  ORIGIN 1.000 0.020 ;
  SIZE 130.695 BY 84.540 ;
  PIN b0
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 23.495 5.200 23.985 5.530 ;
        RECT 2.825 3.280 3.135 3.950 ;
      LAYER met1 ;
        RECT 23.515 5.170 23.965 5.560 ;
        RECT 23.605 5.015 23.895 5.170 ;
        RECT 13.265 4.725 23.895 5.015 ;
        RECT 13.265 4.615 13.555 4.725 ;
        RECT 9.395 4.325 13.555 4.615 ;
        RECT 2.765 3.765 3.195 4.010 ;
        RECT 9.395 3.765 9.685 4.325 ;
        RECT -1.000 3.475 9.685 3.765 ;
        RECT 2.765 3.220 3.195 3.475 ;
    END
  END b0
  PIN b1
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 23.495 13.340 23.985 13.670 ;
        RECT 2.825 11.420 3.135 12.090 ;
      LAYER met1 ;
        RECT 23.515 13.310 23.965 13.700 ;
        RECT 23.605 13.155 23.895 13.310 ;
        RECT 13.265 12.865 23.895 13.155 ;
        RECT 13.265 12.755 13.555 12.865 ;
        RECT 9.395 12.465 13.555 12.755 ;
        RECT 2.765 11.905 3.195 12.150 ;
        RECT 9.395 11.905 9.685 12.465 ;
        RECT -1.000 11.615 9.685 11.905 ;
        RECT 2.765 11.360 3.195 11.615 ;
    END
  END b1
  PIN b2
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 23.495 21.480 23.985 21.810 ;
        RECT 2.825 19.560 3.135 20.230 ;
      LAYER met1 ;
        RECT 23.515 21.450 23.965 21.840 ;
        RECT 23.605 21.295 23.895 21.450 ;
        RECT 13.265 21.005 23.895 21.295 ;
        RECT 13.265 20.895 13.555 21.005 ;
        RECT 9.395 20.605 13.555 20.895 ;
        RECT 2.765 20.045 3.195 20.290 ;
        RECT 9.395 20.045 9.685 20.605 ;
        RECT -1.000 19.755 9.685 20.045 ;
        RECT 2.765 19.500 3.195 19.755 ;
    END
  END b2
  PIN b3
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 23.495 29.620 23.985 29.950 ;
        RECT 2.825 27.700 3.135 28.370 ;
      LAYER met1 ;
        RECT 23.515 29.590 23.965 29.980 ;
        RECT 23.605 29.435 23.895 29.590 ;
        RECT 13.265 29.145 23.895 29.435 ;
        RECT 13.265 29.035 13.555 29.145 ;
        RECT 9.395 28.745 13.555 29.035 ;
        RECT 2.765 28.185 3.195 28.430 ;
        RECT 9.395 28.185 9.685 28.745 ;
        RECT -1.000 27.895 9.685 28.185 ;
        RECT 2.765 27.640 3.195 27.895 ;
    END
  END b3
  PIN b4
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 23.495 37.760 23.985 38.090 ;
        RECT 2.825 35.840 3.135 36.510 ;
      LAYER met1 ;
        RECT 23.515 37.730 23.965 38.120 ;
        RECT 23.605 37.575 23.895 37.730 ;
        RECT 13.265 37.285 23.895 37.575 ;
        RECT 13.265 37.175 13.555 37.285 ;
        RECT 9.395 36.885 13.555 37.175 ;
        RECT 2.765 36.325 3.195 36.570 ;
        RECT 9.395 36.325 9.685 36.885 ;
        RECT -1.000 36.035 9.685 36.325 ;
        RECT 2.765 35.780 3.195 36.035 ;
    END
  END b4
  PIN b5
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 23.495 45.900 23.985 46.230 ;
        RECT 2.825 43.980 3.135 44.650 ;
      LAYER met1 ;
        RECT 23.515 45.870 23.965 46.260 ;
        RECT 23.605 45.715 23.895 45.870 ;
        RECT 13.265 45.425 23.895 45.715 ;
        RECT 13.265 45.315 13.555 45.425 ;
        RECT 9.395 45.025 13.555 45.315 ;
        RECT 2.765 44.465 3.195 44.710 ;
        RECT 9.395 44.465 9.685 45.025 ;
        RECT -1.000 44.175 9.685 44.465 ;
        RECT 2.765 43.920 3.195 44.175 ;
    END
  END b5
  PIN b6
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 23.495 54.040 23.985 54.370 ;
        RECT 2.825 52.120 3.135 52.790 ;
      LAYER met1 ;
        RECT 23.515 54.010 23.965 54.400 ;
        RECT 23.605 53.855 23.895 54.010 ;
        RECT 13.265 53.565 23.895 53.855 ;
        RECT 13.265 53.455 13.555 53.565 ;
        RECT 9.395 53.165 13.555 53.455 ;
        RECT 2.765 52.605 3.195 52.850 ;
        RECT 9.395 52.605 9.685 53.165 ;
        RECT -1.000 52.315 9.685 52.605 ;
        RECT 2.765 52.060 3.195 52.315 ;
    END
  END b6
  PIN b7
    ANTENNAGATEAREA 0.454500 ;
    ANTENNADIFFAREA 0.202500 ;
    PORT
      LAYER li1 ;
        RECT 23.495 62.180 23.985 62.510 ;
        RECT 2.825 60.260 3.135 60.930 ;
      LAYER met1 ;
        RECT 23.515 62.150 23.965 62.540 ;
        RECT 23.605 61.995 23.895 62.150 ;
        RECT 13.265 61.705 23.895 61.995 ;
        RECT 13.265 61.595 13.555 61.705 ;
        RECT 9.395 61.305 13.555 61.595 ;
        RECT 2.765 60.745 3.195 60.990 ;
        RECT 9.395 60.745 9.685 61.305 ;
        RECT -1.000 60.455 9.685 60.745 ;
        RECT 2.765 60.200 3.195 60.455 ;
    END
  END b7
  PIN out
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER li1 ;
        RECT 54.045 68.000 54.215 69.040 ;
        RECT 96.685 68.000 96.855 69.040 ;
        RECT 54.045 66.555 54.215 67.245 ;
        RECT 96.685 66.555 96.855 67.245 ;
      LAYER met1 ;
        RECT 77.180 83.920 78.455 84.520 ;
        RECT 77.380 82.745 78.235 83.920 ;
        RECT 54.015 67.785 54.245 69.020 ;
        RECT 96.655 67.785 96.885 69.020 ;
        RECT 54.000 67.465 54.260 67.785 ;
        RECT 96.640 67.465 96.900 67.785 ;
        RECT 54.015 66.575 54.245 67.465 ;
        RECT 96.655 66.575 96.885 67.465 ;
      LAYER met2 ;
        RECT 77.380 82.745 78.235 83.610 ;
        RECT 53.945 67.485 54.315 67.765 ;
        RECT 96.585 67.485 96.955 67.765 ;
      LAYER met3 ;
        RECT 77.380 82.745 78.235 83.610 ;
        RECT 77.600 77.295 77.900 82.745 ;
        RECT 56.300 76.915 56.620 77.295 ;
        RECT 77.590 76.915 77.910 77.295 ;
        RECT 98.940 76.915 99.260 77.295 ;
        RECT 53.965 67.450 54.295 67.800 ;
        RECT 53.980 66.300 54.280 67.450 ;
        RECT 56.310 66.300 56.610 76.915 ;
        RECT 77.600 76.520 77.900 76.915 ;
        RECT 96.605 67.450 96.935 67.800 ;
        RECT 96.620 66.300 96.920 67.450 ;
        RECT 98.950 66.300 99.250 76.915 ;
        RECT 53.970 65.920 54.290 66.300 ;
        RECT 56.300 65.920 56.620 66.300 ;
        RECT 96.610 65.920 96.930 66.300 ;
        RECT 98.940 65.920 99.260 66.300 ;
      LAYER met4 ;
        RECT 56.295 77.255 56.625 77.270 ;
        RECT 77.585 77.255 77.915 77.270 ;
        RECT 98.935 77.255 99.265 77.270 ;
        RECT 56.295 76.955 99.265 77.255 ;
        RECT 56.295 76.940 56.625 76.955 ;
        RECT 77.585 76.940 77.915 76.955 ;
        RECT 98.935 76.940 99.265 76.955 ;
        RECT 53.965 66.260 54.295 66.275 ;
        RECT 56.295 66.260 56.625 66.275 ;
        RECT 96.605 66.260 96.935 66.275 ;
        RECT 98.935 66.260 99.265 66.275 ;
        RECT 53.525 65.960 56.625 66.260 ;
        RECT 96.165 65.960 99.265 66.260 ;
        RECT 53.965 65.945 54.295 65.960 ;
        RECT 56.295 65.945 56.625 65.960 ;
        RECT 96.605 65.945 96.935 65.960 ;
        RECT 98.935 65.945 99.265 65.960 ;
    END
  END out
  PIN vdd
    ANTENNAGATEAREA 105.000000 ;
    ANTENNADIFFAREA 269.591797 ;
    PORT
      LAYER nwell ;
        RECT 28.730 77.815 129.695 79.390 ;
        RECT 0.000 60.615 1.130 64.985 ;
        RECT 6.665 61.195 22.260 64.985 ;
        RECT 10.130 60.615 22.260 61.195 ;
        RECT 0.000 52.475 1.130 56.845 ;
        RECT 6.665 53.055 22.260 56.845 ;
        RECT 10.130 52.475 22.260 53.055 ;
        RECT 0.000 44.335 1.130 48.705 ;
        RECT 6.665 44.915 22.260 48.705 ;
        RECT 10.130 44.335 22.260 44.915 ;
        RECT 0.000 36.195 1.130 40.565 ;
        RECT 6.665 36.775 22.260 40.565 ;
        RECT 10.130 36.195 22.260 36.775 ;
        RECT 0.000 28.055 1.130 32.425 ;
        RECT 6.665 28.635 22.260 32.425 ;
        RECT 10.130 28.055 22.260 28.635 ;
        RECT 0.000 19.915 1.130 24.285 ;
        RECT 6.665 20.495 22.260 24.285 ;
        RECT 10.130 19.915 22.260 20.495 ;
        RECT 0.000 11.775 1.130 16.145 ;
        RECT 6.665 12.355 22.260 16.145 ;
        RECT 10.130 11.775 22.260 12.355 ;
        RECT 0.000 3.635 1.130 8.005 ;
        RECT 6.665 4.215 22.260 8.005 ;
        RECT 10.130 3.635 22.260 4.215 ;
        RECT 28.730 1.575 30.305 77.815 ;
        RECT 32.325 75.225 35.455 77.815 ;
        RECT 37.650 75.225 40.780 77.815 ;
        RECT 42.985 75.225 46.115 77.815 ;
        RECT 48.310 75.225 51.440 77.815 ;
        RECT 53.645 75.225 56.775 77.815 ;
        RECT 58.970 75.225 62.100 77.815 ;
        RECT 64.305 75.225 67.435 77.815 ;
        RECT 69.630 75.225 72.760 77.815 ;
        RECT 74.965 75.225 78.095 77.815 ;
        RECT 80.290 75.225 83.420 77.815 ;
        RECT 85.625 75.225 88.755 77.815 ;
        RECT 90.950 75.225 94.080 77.815 ;
        RECT 96.285 75.225 99.415 77.815 ;
        RECT 101.610 75.225 104.740 77.815 ;
        RECT 106.945 75.225 110.075 77.815 ;
        RECT 112.270 75.225 115.400 77.815 ;
        RECT 117.605 75.225 120.735 77.815 ;
        RECT 122.930 75.225 126.060 77.815 ;
        RECT 32.335 70.280 35.455 71.905 ;
        RECT 32.325 67.690 35.455 70.280 ;
        RECT 37.660 67.690 40.780 71.905 ;
        RECT 42.995 67.690 46.115 71.905 ;
        RECT 48.320 67.690 51.440 71.905 ;
        RECT 53.655 67.690 56.775 71.905 ;
        RECT 58.980 67.690 62.100 71.905 ;
        RECT 64.315 67.690 67.435 71.905 ;
        RECT 69.640 67.690 72.760 71.905 ;
        RECT 74.975 67.690 78.095 71.905 ;
        RECT 80.300 67.690 83.420 71.905 ;
        RECT 85.635 67.690 88.755 71.905 ;
        RECT 90.960 67.690 94.080 71.905 ;
        RECT 96.295 67.690 99.415 71.905 ;
        RECT 101.620 67.690 104.740 71.905 ;
        RECT 106.955 67.690 110.075 71.905 ;
        RECT 112.280 67.690 115.400 71.905 ;
        RECT 117.615 67.690 120.735 71.905 ;
        RECT 122.940 70.280 126.060 71.905 ;
        RECT 122.930 67.690 126.060 70.280 ;
        RECT 32.335 62.745 35.455 64.370 ;
        RECT 37.660 62.745 40.780 64.370 ;
        RECT 42.995 62.745 46.115 64.370 ;
        RECT 48.320 62.745 51.440 64.370 ;
        RECT 53.655 62.745 56.775 64.370 ;
        RECT 58.980 62.745 62.100 64.370 ;
        RECT 64.315 62.745 67.435 64.370 ;
        RECT 69.640 62.745 72.760 64.370 ;
        RECT 74.975 62.745 78.095 64.370 ;
        RECT 80.300 62.745 83.420 64.370 ;
        RECT 85.635 62.745 88.755 64.370 ;
        RECT 90.960 62.745 94.080 64.370 ;
        RECT 96.295 62.745 99.415 64.370 ;
        RECT 101.620 62.745 104.740 64.370 ;
        RECT 106.955 62.745 110.075 64.370 ;
        RECT 112.280 62.745 115.400 64.370 ;
        RECT 117.615 62.745 120.735 64.370 ;
        RECT 122.940 62.745 126.060 64.370 ;
        RECT 32.325 60.155 35.455 62.745 ;
        RECT 37.650 60.155 40.780 62.745 ;
        RECT 42.985 60.155 46.115 62.745 ;
        RECT 48.310 60.155 51.440 62.745 ;
        RECT 53.645 60.155 56.775 62.745 ;
        RECT 58.970 60.155 62.100 62.745 ;
        RECT 64.305 60.155 67.435 62.745 ;
        RECT 69.630 60.155 72.760 62.745 ;
        RECT 74.965 60.155 78.095 62.745 ;
        RECT 80.290 60.155 83.420 62.745 ;
        RECT 85.625 60.155 88.755 62.745 ;
        RECT 90.950 60.155 94.080 62.745 ;
        RECT 96.285 60.155 99.415 62.745 ;
        RECT 101.610 60.155 104.740 62.745 ;
        RECT 106.945 60.155 110.075 62.745 ;
        RECT 112.270 60.155 115.400 62.745 ;
        RECT 117.605 60.155 120.735 62.745 ;
        RECT 122.930 60.155 126.060 62.745 ;
        RECT 32.335 55.210 35.455 56.835 ;
        RECT 37.660 55.210 40.780 56.835 ;
        RECT 42.995 55.210 46.115 56.835 ;
        RECT 48.320 55.210 51.440 56.835 ;
        RECT 53.655 55.210 56.775 56.835 ;
        RECT 58.980 55.210 62.100 56.835 ;
        RECT 64.315 55.210 67.435 56.835 ;
        RECT 69.640 55.210 72.760 56.835 ;
        RECT 74.975 55.210 78.095 56.835 ;
        RECT 80.300 55.210 83.420 56.835 ;
        RECT 85.635 55.210 88.755 56.835 ;
        RECT 90.960 55.210 94.080 56.835 ;
        RECT 96.295 55.210 99.415 56.835 ;
        RECT 101.620 55.210 104.740 56.835 ;
        RECT 106.955 55.210 110.075 56.835 ;
        RECT 112.280 55.210 115.400 56.835 ;
        RECT 117.615 55.210 120.735 56.835 ;
        RECT 122.940 55.210 126.060 56.835 ;
        RECT 32.325 52.620 35.455 55.210 ;
        RECT 37.650 52.620 40.780 55.210 ;
        RECT 42.985 52.620 46.115 55.210 ;
        RECT 48.310 52.620 51.440 55.210 ;
        RECT 53.645 52.620 56.775 55.210 ;
        RECT 58.970 52.620 62.100 55.210 ;
        RECT 64.305 52.620 67.435 55.210 ;
        RECT 69.630 52.620 72.760 55.210 ;
        RECT 74.965 52.620 78.095 55.210 ;
        RECT 80.290 52.620 83.420 55.210 ;
        RECT 85.625 52.620 88.755 55.210 ;
        RECT 90.950 52.620 94.080 55.210 ;
        RECT 96.285 52.620 99.415 55.210 ;
        RECT 101.610 52.620 104.740 55.210 ;
        RECT 106.945 52.620 110.075 55.210 ;
        RECT 112.270 52.620 115.400 55.210 ;
        RECT 117.605 52.620 120.735 55.210 ;
        RECT 122.930 52.620 126.060 55.210 ;
        RECT 32.335 47.675 35.455 49.300 ;
        RECT 37.660 47.675 40.780 49.300 ;
        RECT 42.995 47.675 46.115 49.300 ;
        RECT 48.320 47.675 51.440 49.300 ;
        RECT 53.655 47.675 56.775 49.300 ;
        RECT 58.980 47.675 62.100 49.300 ;
        RECT 64.315 47.675 67.435 49.300 ;
        RECT 69.640 47.675 72.760 49.300 ;
        RECT 74.975 47.675 78.095 49.300 ;
        RECT 80.300 47.675 83.420 49.300 ;
        RECT 85.635 47.675 88.755 49.300 ;
        RECT 90.960 47.675 94.080 49.300 ;
        RECT 96.295 47.675 99.415 49.300 ;
        RECT 101.620 47.675 104.740 49.300 ;
        RECT 106.955 47.675 110.075 49.300 ;
        RECT 112.280 47.675 115.400 49.300 ;
        RECT 117.615 47.675 120.735 49.300 ;
        RECT 122.940 47.675 126.060 49.300 ;
        RECT 32.325 45.085 35.455 47.675 ;
        RECT 37.650 45.085 40.780 47.675 ;
        RECT 42.985 45.085 46.115 47.675 ;
        RECT 48.310 45.085 51.440 47.675 ;
        RECT 53.645 45.085 56.775 47.675 ;
        RECT 58.970 45.085 62.100 47.675 ;
        RECT 64.305 45.085 67.435 47.675 ;
        RECT 69.630 45.085 72.760 47.675 ;
        RECT 74.965 45.085 78.095 47.675 ;
        RECT 80.290 45.085 83.420 47.675 ;
        RECT 85.625 45.085 88.755 47.675 ;
        RECT 90.950 45.085 94.080 47.675 ;
        RECT 96.285 45.085 99.415 47.675 ;
        RECT 101.610 45.085 104.740 47.675 ;
        RECT 106.945 45.085 110.075 47.675 ;
        RECT 112.270 45.085 115.400 47.675 ;
        RECT 117.605 45.085 120.735 47.675 ;
        RECT 122.930 45.085 126.060 47.675 ;
        RECT 32.335 40.140 35.455 41.765 ;
        RECT 37.660 40.140 40.780 41.765 ;
        RECT 42.995 40.140 46.115 41.765 ;
        RECT 48.320 40.140 51.440 41.765 ;
        RECT 53.655 40.140 56.775 41.765 ;
        RECT 58.980 40.140 62.100 41.765 ;
        RECT 64.315 40.140 67.435 41.765 ;
        RECT 69.640 40.140 72.760 41.765 ;
        RECT 74.975 40.140 78.095 41.765 ;
        RECT 80.300 40.140 83.420 41.765 ;
        RECT 85.635 40.140 88.755 41.765 ;
        RECT 90.960 40.140 94.080 41.765 ;
        RECT 96.295 40.140 99.415 41.765 ;
        RECT 101.620 40.140 104.740 41.765 ;
        RECT 106.955 40.140 110.075 41.765 ;
        RECT 112.280 40.140 115.400 41.765 ;
        RECT 117.615 40.140 120.735 41.765 ;
        RECT 122.940 40.140 126.060 41.765 ;
        RECT 32.325 37.550 35.455 40.140 ;
        RECT 37.650 37.550 40.780 40.140 ;
        RECT 42.985 37.550 46.115 40.140 ;
        RECT 48.310 37.550 51.440 40.140 ;
        RECT 53.645 37.550 56.775 40.140 ;
        RECT 58.970 37.550 62.100 40.140 ;
        RECT 64.305 37.550 67.435 40.140 ;
        RECT 69.630 37.550 72.760 40.140 ;
        RECT 74.965 37.550 78.095 40.140 ;
        RECT 80.290 37.550 83.420 40.140 ;
        RECT 85.625 37.550 88.755 40.140 ;
        RECT 90.950 37.550 94.080 40.140 ;
        RECT 96.285 37.550 99.415 40.140 ;
        RECT 101.610 37.550 104.740 40.140 ;
        RECT 106.945 37.550 110.075 40.140 ;
        RECT 112.270 37.550 115.400 40.140 ;
        RECT 117.605 37.550 120.735 40.140 ;
        RECT 122.930 37.550 126.060 40.140 ;
        RECT 32.335 32.605 35.455 34.230 ;
        RECT 37.660 32.605 40.780 34.230 ;
        RECT 42.995 32.605 46.115 34.230 ;
        RECT 48.320 32.605 51.440 34.230 ;
        RECT 53.655 32.605 56.775 34.230 ;
        RECT 58.980 32.605 62.100 34.230 ;
        RECT 64.315 32.605 67.435 34.230 ;
        RECT 69.640 32.605 72.760 34.230 ;
        RECT 74.975 32.605 78.095 34.230 ;
        RECT 80.300 32.605 83.420 34.230 ;
        RECT 85.635 32.605 88.755 34.230 ;
        RECT 90.960 32.605 94.080 34.230 ;
        RECT 96.295 32.605 99.415 34.230 ;
        RECT 101.620 32.605 104.740 34.230 ;
        RECT 106.955 32.605 110.075 34.230 ;
        RECT 112.280 32.605 115.400 34.230 ;
        RECT 117.615 32.605 120.735 34.230 ;
        RECT 122.940 32.605 126.060 34.230 ;
        RECT 32.325 30.015 35.455 32.605 ;
        RECT 37.650 30.015 40.780 32.605 ;
        RECT 42.985 30.015 46.115 32.605 ;
        RECT 48.310 30.015 51.440 32.605 ;
        RECT 53.645 30.015 56.775 32.605 ;
        RECT 58.970 30.015 62.100 32.605 ;
        RECT 64.305 30.015 67.435 32.605 ;
        RECT 69.630 30.015 72.760 32.605 ;
        RECT 74.965 30.015 78.095 32.605 ;
        RECT 80.290 30.015 83.420 32.605 ;
        RECT 85.625 30.015 88.755 32.605 ;
        RECT 90.950 30.015 94.080 32.605 ;
        RECT 96.285 30.015 99.415 32.605 ;
        RECT 101.610 30.015 104.740 32.605 ;
        RECT 106.945 30.015 110.075 32.605 ;
        RECT 112.270 30.015 115.400 32.605 ;
        RECT 117.605 30.015 120.735 32.605 ;
        RECT 122.930 30.015 126.060 32.605 ;
        RECT 32.335 25.070 35.455 26.695 ;
        RECT 37.660 25.070 40.780 26.695 ;
        RECT 42.995 25.070 46.115 26.695 ;
        RECT 48.320 25.070 51.440 26.695 ;
        RECT 53.655 25.070 56.775 26.695 ;
        RECT 58.980 25.070 62.100 26.695 ;
        RECT 64.315 25.070 67.435 26.695 ;
        RECT 69.640 25.070 72.760 26.695 ;
        RECT 74.975 25.070 78.095 26.695 ;
        RECT 80.300 25.070 83.420 26.695 ;
        RECT 85.635 25.070 88.755 26.695 ;
        RECT 90.960 25.070 94.080 26.695 ;
        RECT 96.295 25.070 99.415 26.695 ;
        RECT 101.620 25.070 104.740 26.695 ;
        RECT 106.955 25.070 110.075 26.695 ;
        RECT 112.280 25.070 115.400 26.695 ;
        RECT 117.615 25.070 120.735 26.695 ;
        RECT 122.940 25.070 126.060 26.695 ;
        RECT 32.325 22.480 35.455 25.070 ;
        RECT 37.650 22.480 40.780 25.070 ;
        RECT 42.985 22.480 46.115 25.070 ;
        RECT 48.310 22.480 51.440 25.070 ;
        RECT 53.645 22.480 56.775 25.070 ;
        RECT 58.970 22.480 62.100 25.070 ;
        RECT 64.305 22.480 67.435 25.070 ;
        RECT 69.630 22.480 72.760 25.070 ;
        RECT 74.965 22.480 78.095 25.070 ;
        RECT 80.290 22.480 83.420 25.070 ;
        RECT 85.625 22.480 88.755 25.070 ;
        RECT 90.950 22.480 94.080 25.070 ;
        RECT 96.285 22.480 99.415 25.070 ;
        RECT 101.610 22.480 104.740 25.070 ;
        RECT 106.945 22.480 110.075 25.070 ;
        RECT 112.270 22.480 115.400 25.070 ;
        RECT 117.605 22.480 120.735 25.070 ;
        RECT 122.930 22.480 126.060 25.070 ;
        RECT 32.335 17.535 35.455 19.160 ;
        RECT 37.660 17.535 40.780 19.160 ;
        RECT 32.325 14.945 35.455 17.535 ;
        RECT 37.650 14.945 40.780 17.535 ;
        RECT 42.995 15.785 46.115 19.160 ;
        RECT 48.320 17.535 51.440 19.160 ;
        RECT 42.985 14.945 46.115 15.785 ;
        RECT 48.310 14.945 51.440 17.535 ;
        RECT 53.655 15.785 56.775 19.160 ;
        RECT 58.980 17.535 62.100 19.160 ;
        RECT 53.645 14.945 56.775 15.785 ;
        RECT 58.970 14.945 62.100 17.535 ;
        RECT 64.315 15.785 67.435 19.160 ;
        RECT 69.640 17.535 72.760 19.160 ;
        RECT 64.305 14.945 67.435 15.785 ;
        RECT 69.630 14.945 72.760 17.535 ;
        RECT 74.975 15.785 78.095 19.160 ;
        RECT 80.300 17.535 83.420 19.160 ;
        RECT 74.965 14.945 78.095 15.785 ;
        RECT 80.290 14.945 83.420 17.535 ;
        RECT 85.635 15.785 88.755 19.160 ;
        RECT 90.960 17.535 94.080 19.160 ;
        RECT 85.625 14.945 88.755 15.785 ;
        RECT 90.950 14.945 94.080 17.535 ;
        RECT 96.295 15.785 99.415 19.160 ;
        RECT 101.620 17.535 104.740 19.160 ;
        RECT 96.285 14.945 99.415 15.785 ;
        RECT 101.610 14.945 104.740 17.535 ;
        RECT 106.955 15.785 110.075 19.160 ;
        RECT 112.280 17.535 115.400 19.160 ;
        RECT 106.945 14.945 110.075 15.785 ;
        RECT 112.270 14.945 115.400 17.535 ;
        RECT 117.615 15.785 120.735 19.160 ;
        RECT 122.940 17.535 126.060 19.160 ;
        RECT 117.605 14.945 120.735 15.785 ;
        RECT 122.930 14.945 126.060 17.535 ;
        RECT 32.335 10.000 35.455 11.625 ;
        RECT 37.660 10.000 40.780 11.625 ;
        RECT 42.995 10.000 46.115 11.625 ;
        RECT 48.320 10.000 51.440 11.625 ;
        RECT 53.655 10.000 56.775 11.625 ;
        RECT 58.980 10.000 62.100 11.625 ;
        RECT 64.315 10.000 67.435 11.625 ;
        RECT 69.640 10.000 72.760 11.625 ;
        RECT 74.975 10.000 78.095 11.625 ;
        RECT 80.300 10.000 83.420 11.625 ;
        RECT 85.635 10.000 88.755 11.625 ;
        RECT 90.960 10.000 94.080 11.625 ;
        RECT 96.295 10.000 99.415 11.625 ;
        RECT 101.620 10.000 104.740 11.625 ;
        RECT 106.955 10.000 110.075 11.625 ;
        RECT 112.280 10.000 115.400 11.625 ;
        RECT 117.615 10.000 120.735 11.625 ;
        RECT 122.940 10.000 126.060 11.625 ;
        RECT 32.325 7.410 35.455 10.000 ;
        RECT 37.650 7.410 40.780 10.000 ;
        RECT 42.985 7.410 46.115 10.000 ;
        RECT 48.310 7.410 51.440 10.000 ;
        RECT 53.645 7.410 56.775 10.000 ;
        RECT 58.970 7.410 62.100 10.000 ;
        RECT 64.305 7.410 67.435 10.000 ;
        RECT 69.630 7.410 72.760 10.000 ;
        RECT 74.965 7.410 78.095 10.000 ;
        RECT 80.290 7.410 83.420 10.000 ;
        RECT 85.625 7.410 88.755 10.000 ;
        RECT 90.950 7.410 94.080 10.000 ;
        RECT 96.285 7.410 99.415 10.000 ;
        RECT 101.610 7.410 104.740 10.000 ;
        RECT 106.945 7.410 110.075 10.000 ;
        RECT 112.270 7.410 115.400 10.000 ;
        RECT 117.605 7.410 120.735 10.000 ;
        RECT 122.930 7.410 126.060 10.000 ;
        RECT 32.335 1.575 35.455 4.090 ;
        RECT 37.660 1.575 40.780 4.090 ;
        RECT 42.995 1.575 46.115 4.090 ;
        RECT 48.320 1.575 51.440 4.090 ;
        RECT 53.655 1.575 56.775 4.090 ;
        RECT 58.980 1.575 62.100 4.090 ;
        RECT 64.315 1.575 67.435 4.090 ;
        RECT 69.640 1.575 72.760 4.090 ;
        RECT 74.975 1.575 78.095 4.090 ;
        RECT 80.300 1.575 83.420 4.090 ;
        RECT 85.635 1.575 88.755 4.090 ;
        RECT 90.960 1.575 94.080 4.090 ;
        RECT 96.295 1.575 99.415 4.090 ;
        RECT 101.620 1.575 104.740 4.090 ;
        RECT 106.955 1.575 110.075 4.090 ;
        RECT 112.280 1.575 115.400 4.090 ;
        RECT 117.615 1.575 120.735 4.090 ;
        RECT 122.940 1.575 126.060 4.090 ;
        RECT 128.120 1.575 129.695 77.815 ;
        RECT 28.730 0.000 129.695 1.575 ;
      LAYER li1 ;
        RECT 29.160 78.790 129.265 78.960 ;
        RECT 8.085 63.135 8.675 63.530 ;
        RECT 9.540 63.135 10.130 64.675 ;
        RECT 10.980 63.115 11.570 64.695 ;
        RECT 12.440 63.115 13.390 64.590 ;
        RECT 14.010 63.115 14.600 64.590 ;
        RECT 14.825 63.245 15.715 64.425 ;
        RECT 16.505 63.245 17.395 64.485 ;
        RECT 18.065 63.245 18.955 64.485 ;
        RECT 19.625 63.245 20.515 64.485 ;
        RECT 21.185 63.245 21.755 64.485 ;
        RECT 14.825 63.075 21.755 63.245 ;
        RECT 0.330 62.715 1.130 62.885 ;
        RECT 8.085 62.715 21.930 62.885 ;
        RECT 8.335 61.525 8.925 62.435 ;
        RECT 11.000 60.905 11.950 62.485 ;
        RECT 12.570 60.905 13.160 62.485 ;
        RECT 13.385 62.355 20.315 62.525 ;
        RECT 13.385 61.175 14.275 62.355 ;
        RECT 15.065 61.115 15.955 62.355 ;
        RECT 16.625 61.115 17.515 62.355 ;
        RECT 18.185 61.115 19.075 62.355 ;
        RECT 19.745 61.115 20.315 62.355 ;
        RECT 8.085 54.995 8.675 55.390 ;
        RECT 9.540 54.995 10.130 56.535 ;
        RECT 10.980 54.975 11.570 56.555 ;
        RECT 12.440 54.975 13.390 56.450 ;
        RECT 14.010 54.975 14.600 56.450 ;
        RECT 14.825 55.105 15.715 56.285 ;
        RECT 16.505 55.105 17.395 56.345 ;
        RECT 18.065 55.105 18.955 56.345 ;
        RECT 19.625 55.105 20.515 56.345 ;
        RECT 21.185 55.105 21.755 56.345 ;
        RECT 14.825 54.935 21.755 55.105 ;
        RECT 0.330 54.575 1.130 54.745 ;
        RECT 8.085 54.575 21.930 54.745 ;
        RECT 8.335 53.385 8.925 54.295 ;
        RECT 11.000 52.765 11.950 54.345 ;
        RECT 12.570 52.765 13.160 54.345 ;
        RECT 13.385 54.215 20.315 54.385 ;
        RECT 13.385 53.035 14.275 54.215 ;
        RECT 15.065 52.975 15.955 54.215 ;
        RECT 16.625 52.975 17.515 54.215 ;
        RECT 18.185 52.975 19.075 54.215 ;
        RECT 19.745 52.975 20.315 54.215 ;
        RECT 8.085 46.855 8.675 47.250 ;
        RECT 9.540 46.855 10.130 48.395 ;
        RECT 10.980 46.835 11.570 48.415 ;
        RECT 12.440 46.835 13.390 48.310 ;
        RECT 14.010 46.835 14.600 48.310 ;
        RECT 14.825 46.965 15.715 48.145 ;
        RECT 16.505 46.965 17.395 48.205 ;
        RECT 18.065 46.965 18.955 48.205 ;
        RECT 19.625 46.965 20.515 48.205 ;
        RECT 21.185 46.965 21.755 48.205 ;
        RECT 14.825 46.795 21.755 46.965 ;
        RECT 0.330 46.435 1.130 46.605 ;
        RECT 8.085 46.435 21.930 46.605 ;
        RECT 8.335 45.245 8.925 46.155 ;
        RECT 11.000 44.625 11.950 46.205 ;
        RECT 12.570 44.625 13.160 46.205 ;
        RECT 13.385 46.075 20.315 46.245 ;
        RECT 13.385 44.895 14.275 46.075 ;
        RECT 15.065 44.835 15.955 46.075 ;
        RECT 16.625 44.835 17.515 46.075 ;
        RECT 18.185 44.835 19.075 46.075 ;
        RECT 19.745 44.835 20.315 46.075 ;
        RECT 8.085 38.715 8.675 39.110 ;
        RECT 9.540 38.715 10.130 40.255 ;
        RECT 10.980 38.695 11.570 40.275 ;
        RECT 12.440 38.695 13.390 40.170 ;
        RECT 14.010 38.695 14.600 40.170 ;
        RECT 14.825 38.825 15.715 40.005 ;
        RECT 16.505 38.825 17.395 40.065 ;
        RECT 18.065 38.825 18.955 40.065 ;
        RECT 19.625 38.825 20.515 40.065 ;
        RECT 21.185 38.825 21.755 40.065 ;
        RECT 14.825 38.655 21.755 38.825 ;
        RECT 0.330 38.295 1.130 38.465 ;
        RECT 8.085 38.295 21.930 38.465 ;
        RECT 8.335 37.105 8.925 38.015 ;
        RECT 11.000 36.485 11.950 38.065 ;
        RECT 12.570 36.485 13.160 38.065 ;
        RECT 13.385 37.935 20.315 38.105 ;
        RECT 13.385 36.755 14.275 37.935 ;
        RECT 15.065 36.695 15.955 37.935 ;
        RECT 16.625 36.695 17.515 37.935 ;
        RECT 18.185 36.695 19.075 37.935 ;
        RECT 19.745 36.695 20.315 37.935 ;
        RECT 8.085 30.575 8.675 30.970 ;
        RECT 9.540 30.575 10.130 32.115 ;
        RECT 10.980 30.555 11.570 32.135 ;
        RECT 12.440 30.555 13.390 32.030 ;
        RECT 14.010 30.555 14.600 32.030 ;
        RECT 14.825 30.685 15.715 31.865 ;
        RECT 16.505 30.685 17.395 31.925 ;
        RECT 18.065 30.685 18.955 31.925 ;
        RECT 19.625 30.685 20.515 31.925 ;
        RECT 21.185 30.685 21.755 31.925 ;
        RECT 14.825 30.515 21.755 30.685 ;
        RECT 0.330 30.155 1.130 30.325 ;
        RECT 8.085 30.155 21.930 30.325 ;
        RECT 8.335 28.965 8.925 29.875 ;
        RECT 11.000 28.345 11.950 29.925 ;
        RECT 12.570 28.345 13.160 29.925 ;
        RECT 13.385 29.795 20.315 29.965 ;
        RECT 13.385 28.615 14.275 29.795 ;
        RECT 15.065 28.555 15.955 29.795 ;
        RECT 16.625 28.555 17.515 29.795 ;
        RECT 18.185 28.555 19.075 29.795 ;
        RECT 19.745 28.555 20.315 29.795 ;
        RECT 8.085 22.435 8.675 22.830 ;
        RECT 9.540 22.435 10.130 23.975 ;
        RECT 10.980 22.415 11.570 23.995 ;
        RECT 12.440 22.415 13.390 23.890 ;
        RECT 14.010 22.415 14.600 23.890 ;
        RECT 14.825 22.545 15.715 23.725 ;
        RECT 16.505 22.545 17.395 23.785 ;
        RECT 18.065 22.545 18.955 23.785 ;
        RECT 19.625 22.545 20.515 23.785 ;
        RECT 21.185 22.545 21.755 23.785 ;
        RECT 14.825 22.375 21.755 22.545 ;
        RECT 0.330 22.015 1.130 22.185 ;
        RECT 8.085 22.015 21.930 22.185 ;
        RECT 8.335 20.825 8.925 21.735 ;
        RECT 11.000 20.205 11.950 21.785 ;
        RECT 12.570 20.205 13.160 21.785 ;
        RECT 13.385 21.655 20.315 21.825 ;
        RECT 13.385 20.475 14.275 21.655 ;
        RECT 15.065 20.415 15.955 21.655 ;
        RECT 16.625 20.415 17.515 21.655 ;
        RECT 18.185 20.415 19.075 21.655 ;
        RECT 19.745 20.415 20.315 21.655 ;
        RECT 8.085 14.295 8.675 14.690 ;
        RECT 9.540 14.295 10.130 15.835 ;
        RECT 10.980 14.275 11.570 15.855 ;
        RECT 12.440 14.275 13.390 15.750 ;
        RECT 14.010 14.275 14.600 15.750 ;
        RECT 14.825 14.405 15.715 15.585 ;
        RECT 16.505 14.405 17.395 15.645 ;
        RECT 18.065 14.405 18.955 15.645 ;
        RECT 19.625 14.405 20.515 15.645 ;
        RECT 21.185 14.405 21.755 15.645 ;
        RECT 14.825 14.235 21.755 14.405 ;
        RECT 0.330 13.875 1.130 14.045 ;
        RECT 8.085 13.875 21.930 14.045 ;
        RECT 8.335 12.685 8.925 13.595 ;
        RECT 11.000 12.065 11.950 13.645 ;
        RECT 12.570 12.065 13.160 13.645 ;
        RECT 13.385 13.515 20.315 13.685 ;
        RECT 13.385 12.335 14.275 13.515 ;
        RECT 15.065 12.275 15.955 13.515 ;
        RECT 16.625 12.275 17.515 13.515 ;
        RECT 18.185 12.275 19.075 13.515 ;
        RECT 19.745 12.275 20.315 13.515 ;
        RECT 8.085 6.155 8.675 6.550 ;
        RECT 9.540 6.155 10.130 7.695 ;
        RECT 10.980 6.135 11.570 7.715 ;
        RECT 12.440 6.135 13.390 7.610 ;
        RECT 14.010 6.135 14.600 7.610 ;
        RECT 14.825 6.265 15.715 7.445 ;
        RECT 16.505 6.265 17.395 7.505 ;
        RECT 18.065 6.265 18.955 7.505 ;
        RECT 19.625 6.265 20.515 7.505 ;
        RECT 21.185 6.265 21.755 7.505 ;
        RECT 14.825 6.095 21.755 6.265 ;
        RECT 0.330 5.735 1.130 5.905 ;
        RECT 8.085 5.735 21.930 5.905 ;
        RECT 8.335 4.545 8.925 5.455 ;
        RECT 11.000 3.925 11.950 5.505 ;
        RECT 12.570 3.925 13.160 5.505 ;
        RECT 13.385 5.375 20.315 5.545 ;
        RECT 13.385 4.195 14.275 5.375 ;
        RECT 15.065 4.135 15.955 5.375 ;
        RECT 16.625 4.135 17.515 5.375 ;
        RECT 18.185 4.135 19.075 5.375 ;
        RECT 19.745 4.135 20.315 5.375 ;
        RECT 29.160 0.600 29.330 78.790 ;
        RECT 33.225 77.255 34.580 77.485 ;
        RECT 38.550 77.255 39.905 77.485 ;
        RECT 43.885 77.255 45.240 77.485 ;
        RECT 49.210 77.255 50.565 77.485 ;
        RECT 54.545 77.255 55.900 77.485 ;
        RECT 59.870 77.255 61.225 77.485 ;
        RECT 65.205 77.255 66.560 77.485 ;
        RECT 70.530 77.255 71.885 77.485 ;
        RECT 75.865 77.255 77.220 77.485 ;
        RECT 81.190 77.255 82.545 77.485 ;
        RECT 86.525 77.255 87.880 77.485 ;
        RECT 91.850 77.255 93.205 77.485 ;
        RECT 97.185 77.255 98.540 77.485 ;
        RECT 102.510 77.255 103.865 77.485 ;
        RECT 107.845 77.255 109.200 77.485 ;
        RECT 113.170 77.255 114.525 77.485 ;
        RECT 118.505 77.255 119.860 77.485 ;
        RECT 123.830 77.255 125.185 77.485 ;
        RECT 32.955 76.790 33.455 76.960 ;
        RECT 33.810 76.875 34.005 77.255 ;
        RECT 34.335 76.790 34.835 76.960 ;
        RECT 38.280 76.790 38.780 76.960 ;
        RECT 39.135 76.875 39.330 77.255 ;
        RECT 39.660 76.790 40.160 76.960 ;
        RECT 43.615 76.790 44.115 76.960 ;
        RECT 44.470 76.875 44.665 77.255 ;
        RECT 44.995 76.790 45.495 76.960 ;
        RECT 48.940 76.790 49.440 76.960 ;
        RECT 49.795 76.875 49.990 77.255 ;
        RECT 50.320 76.790 50.820 76.960 ;
        RECT 54.275 76.790 54.775 76.960 ;
        RECT 55.130 76.875 55.325 77.255 ;
        RECT 55.655 76.790 56.155 76.960 ;
        RECT 59.600 76.790 60.100 76.960 ;
        RECT 60.455 76.875 60.650 77.255 ;
        RECT 60.980 76.790 61.480 76.960 ;
        RECT 64.935 76.790 65.435 76.960 ;
        RECT 65.790 76.875 65.985 77.255 ;
        RECT 66.315 76.790 66.815 76.960 ;
        RECT 70.260 76.790 70.760 76.960 ;
        RECT 71.115 76.875 71.310 77.255 ;
        RECT 71.640 76.790 72.140 76.960 ;
        RECT 75.595 76.790 76.095 76.960 ;
        RECT 76.450 76.875 76.645 77.255 ;
        RECT 76.975 76.790 77.475 76.960 ;
        RECT 80.920 76.790 81.420 76.960 ;
        RECT 81.775 76.875 81.970 77.255 ;
        RECT 82.300 76.790 82.800 76.960 ;
        RECT 86.255 76.790 86.755 76.960 ;
        RECT 87.110 76.875 87.305 77.255 ;
        RECT 87.635 76.790 88.135 76.960 ;
        RECT 91.580 76.790 92.080 76.960 ;
        RECT 92.435 76.875 92.630 77.255 ;
        RECT 92.960 76.790 93.460 76.960 ;
        RECT 96.915 76.790 97.415 76.960 ;
        RECT 97.770 76.875 97.965 77.255 ;
        RECT 98.295 76.790 98.795 76.960 ;
        RECT 102.240 76.790 102.740 76.960 ;
        RECT 103.095 76.875 103.290 77.255 ;
        RECT 103.620 76.790 104.120 76.960 ;
        RECT 107.575 76.790 108.075 76.960 ;
        RECT 108.430 76.875 108.625 77.255 ;
        RECT 108.955 76.790 109.455 76.960 ;
        RECT 112.900 76.790 113.400 76.960 ;
        RECT 113.755 76.875 113.950 77.255 ;
        RECT 114.280 76.790 114.780 76.960 ;
        RECT 118.235 76.790 118.735 76.960 ;
        RECT 119.090 76.875 119.285 77.255 ;
        RECT 119.615 76.790 120.115 76.960 ;
        RECT 123.560 76.790 124.060 76.960 ;
        RECT 124.415 76.875 124.610 77.255 ;
        RECT 124.940 76.790 125.440 76.960 ;
        RECT 32.955 70.170 33.455 70.340 ;
        RECT 33.810 69.950 34.005 70.340 ;
        RECT 34.335 70.170 34.835 70.340 ;
        RECT 38.280 70.170 38.780 70.340 ;
        RECT 39.135 69.950 39.330 70.340 ;
        RECT 39.660 70.170 40.160 70.340 ;
        RECT 43.615 70.170 44.115 70.340 ;
        RECT 44.470 69.950 44.665 70.340 ;
        RECT 44.995 70.170 45.495 70.340 ;
        RECT 48.940 70.170 49.440 70.340 ;
        RECT 49.795 69.950 49.990 70.340 ;
        RECT 50.320 70.170 50.820 70.340 ;
        RECT 54.275 70.170 54.775 70.340 ;
        RECT 55.130 69.950 55.325 70.340 ;
        RECT 55.655 70.170 56.155 70.340 ;
        RECT 59.600 70.170 60.100 70.340 ;
        RECT 60.455 69.950 60.650 70.340 ;
        RECT 60.980 70.170 61.480 70.340 ;
        RECT 64.935 70.170 65.435 70.340 ;
        RECT 65.790 69.950 65.985 70.340 ;
        RECT 66.315 70.170 66.815 70.340 ;
        RECT 70.260 70.170 70.760 70.340 ;
        RECT 71.115 69.950 71.310 70.340 ;
        RECT 71.640 70.170 72.140 70.340 ;
        RECT 75.595 70.170 76.095 70.340 ;
        RECT 76.450 69.950 76.645 70.340 ;
        RECT 76.975 70.170 77.475 70.340 ;
        RECT 80.920 70.170 81.420 70.340 ;
        RECT 81.775 69.950 81.970 70.340 ;
        RECT 82.300 70.170 82.800 70.340 ;
        RECT 86.255 70.170 86.755 70.340 ;
        RECT 87.110 69.950 87.305 70.340 ;
        RECT 87.635 70.170 88.135 70.340 ;
        RECT 91.580 70.170 92.080 70.340 ;
        RECT 92.435 69.950 92.630 70.340 ;
        RECT 92.960 70.170 93.460 70.340 ;
        RECT 96.915 70.170 97.415 70.340 ;
        RECT 97.770 69.950 97.965 70.340 ;
        RECT 98.295 70.170 98.795 70.340 ;
        RECT 102.240 70.170 102.740 70.340 ;
        RECT 103.095 69.950 103.290 70.340 ;
        RECT 103.620 70.170 104.120 70.340 ;
        RECT 107.575 70.170 108.075 70.340 ;
        RECT 108.430 69.950 108.625 70.340 ;
        RECT 108.955 70.170 109.455 70.340 ;
        RECT 112.900 70.170 113.400 70.340 ;
        RECT 113.755 69.950 113.950 70.340 ;
        RECT 114.280 70.170 114.780 70.340 ;
        RECT 118.235 70.170 118.735 70.340 ;
        RECT 119.090 69.950 119.285 70.340 ;
        RECT 119.615 70.170 120.115 70.340 ;
        RECT 123.560 70.170 124.060 70.340 ;
        RECT 124.415 69.950 124.610 70.340 ;
        RECT 124.940 70.170 125.440 70.340 ;
        RECT 33.225 69.720 34.580 69.950 ;
        RECT 38.550 69.720 39.905 69.950 ;
        RECT 43.885 69.720 45.240 69.950 ;
        RECT 49.210 69.720 50.565 69.950 ;
        RECT 54.545 69.720 55.900 69.950 ;
        RECT 59.870 69.720 61.225 69.950 ;
        RECT 65.205 69.720 66.560 69.950 ;
        RECT 70.530 69.720 71.885 69.950 ;
        RECT 75.865 69.720 77.220 69.950 ;
        RECT 81.190 69.720 82.545 69.950 ;
        RECT 86.525 69.720 87.880 69.950 ;
        RECT 91.850 69.720 93.205 69.950 ;
        RECT 97.185 69.720 98.540 69.950 ;
        RECT 102.510 69.720 103.865 69.950 ;
        RECT 107.845 69.720 109.200 69.950 ;
        RECT 113.170 69.720 114.525 69.950 ;
        RECT 118.505 69.720 119.860 69.950 ;
        RECT 123.830 69.720 125.185 69.950 ;
        RECT 32.955 69.255 33.455 69.425 ;
        RECT 33.810 69.340 34.005 69.720 ;
        RECT 34.335 69.255 34.835 69.425 ;
        RECT 39.135 69.340 39.330 69.720 ;
        RECT 44.470 69.340 44.665 69.720 ;
        RECT 49.795 69.340 49.990 69.720 ;
        RECT 55.130 69.340 55.325 69.720 ;
        RECT 60.455 69.340 60.650 69.720 ;
        RECT 65.790 69.340 65.985 69.720 ;
        RECT 71.115 69.340 71.310 69.720 ;
        RECT 75.595 69.255 76.095 69.425 ;
        RECT 76.450 69.340 76.645 69.720 ;
        RECT 81.775 69.340 81.970 69.720 ;
        RECT 87.110 69.340 87.305 69.720 ;
        RECT 92.435 69.340 92.630 69.720 ;
        RECT 97.770 69.340 97.965 69.720 ;
        RECT 103.095 69.340 103.290 69.720 ;
        RECT 108.430 69.340 108.625 69.720 ;
        RECT 113.755 69.340 113.950 69.720 ;
        RECT 118.235 69.255 118.735 69.425 ;
        RECT 119.090 69.340 119.285 69.720 ;
        RECT 123.560 69.255 124.060 69.425 ;
        RECT 124.415 69.340 124.610 69.720 ;
        RECT 124.940 69.255 125.440 69.425 ;
        RECT 32.955 62.635 33.455 62.805 ;
        RECT 33.810 62.415 34.005 62.805 ;
        RECT 34.335 62.635 34.835 62.805 ;
        RECT 39.135 62.415 39.330 62.805 ;
        RECT 44.470 62.415 44.665 62.805 ;
        RECT 49.795 62.415 49.990 62.805 ;
        RECT 55.130 62.415 55.325 62.805 ;
        RECT 60.455 62.415 60.650 62.805 ;
        RECT 65.790 62.415 65.985 62.805 ;
        RECT 71.115 62.415 71.310 62.805 ;
        RECT 76.450 62.415 76.645 62.805 ;
        RECT 81.775 62.415 81.970 62.805 ;
        RECT 87.110 62.415 87.305 62.805 ;
        RECT 92.435 62.415 92.630 62.805 ;
        RECT 97.770 62.415 97.965 62.805 ;
        RECT 103.095 62.415 103.290 62.805 ;
        RECT 108.430 62.415 108.625 62.805 ;
        RECT 113.755 62.415 113.950 62.805 ;
        RECT 119.090 62.415 119.285 62.805 ;
        RECT 123.560 62.635 124.060 62.805 ;
        RECT 124.415 62.415 124.610 62.805 ;
        RECT 124.940 62.635 125.440 62.805 ;
        RECT 33.225 62.185 34.580 62.415 ;
        RECT 38.550 62.185 39.905 62.415 ;
        RECT 43.885 62.185 45.240 62.415 ;
        RECT 49.210 62.185 50.565 62.415 ;
        RECT 54.545 62.185 55.900 62.415 ;
        RECT 59.870 62.185 61.225 62.415 ;
        RECT 65.205 62.185 66.560 62.415 ;
        RECT 70.530 62.185 71.885 62.415 ;
        RECT 75.865 62.185 77.220 62.415 ;
        RECT 81.190 62.185 82.545 62.415 ;
        RECT 86.525 62.185 87.880 62.415 ;
        RECT 91.850 62.185 93.205 62.415 ;
        RECT 97.185 62.185 98.540 62.415 ;
        RECT 102.510 62.185 103.865 62.415 ;
        RECT 107.845 62.185 109.200 62.415 ;
        RECT 113.170 62.185 114.525 62.415 ;
        RECT 118.505 62.185 119.860 62.415 ;
        RECT 123.830 62.185 125.185 62.415 ;
        RECT 32.955 61.720 33.455 61.890 ;
        RECT 33.810 61.805 34.005 62.185 ;
        RECT 34.335 61.720 34.835 61.890 ;
        RECT 39.135 61.805 39.330 62.185 ;
        RECT 44.470 61.805 44.665 62.185 ;
        RECT 49.795 61.805 49.990 62.185 ;
        RECT 55.130 61.805 55.325 62.185 ;
        RECT 60.455 61.805 60.650 62.185 ;
        RECT 65.790 61.805 65.985 62.185 ;
        RECT 71.115 61.805 71.310 62.185 ;
        RECT 76.450 61.805 76.645 62.185 ;
        RECT 81.775 61.805 81.970 62.185 ;
        RECT 87.110 61.805 87.305 62.185 ;
        RECT 92.435 61.805 92.630 62.185 ;
        RECT 97.770 61.805 97.965 62.185 ;
        RECT 103.095 61.805 103.290 62.185 ;
        RECT 108.430 61.805 108.625 62.185 ;
        RECT 113.755 61.805 113.950 62.185 ;
        RECT 119.090 61.805 119.285 62.185 ;
        RECT 123.560 61.720 124.060 61.890 ;
        RECT 124.415 61.805 124.610 62.185 ;
        RECT 124.940 61.720 125.440 61.890 ;
        RECT 32.955 55.100 33.455 55.270 ;
        RECT 33.810 54.880 34.005 55.270 ;
        RECT 34.335 55.100 34.835 55.270 ;
        RECT 39.135 54.880 39.330 55.270 ;
        RECT 44.470 54.880 44.665 55.270 ;
        RECT 49.795 54.880 49.990 55.270 ;
        RECT 55.130 54.880 55.325 55.270 ;
        RECT 60.455 54.880 60.650 55.270 ;
        RECT 65.790 54.880 65.985 55.270 ;
        RECT 71.115 54.880 71.310 55.270 ;
        RECT 76.450 54.880 76.645 55.270 ;
        RECT 81.775 54.880 81.970 55.270 ;
        RECT 87.110 54.880 87.305 55.270 ;
        RECT 92.435 54.880 92.630 55.270 ;
        RECT 97.770 54.880 97.965 55.270 ;
        RECT 103.095 54.880 103.290 55.270 ;
        RECT 108.430 54.880 108.625 55.270 ;
        RECT 113.755 54.880 113.950 55.270 ;
        RECT 119.090 54.880 119.285 55.270 ;
        RECT 123.560 55.100 124.060 55.270 ;
        RECT 124.415 54.880 124.610 55.270 ;
        RECT 124.940 55.100 125.440 55.270 ;
        RECT 33.225 54.650 34.580 54.880 ;
        RECT 38.550 54.650 39.905 54.880 ;
        RECT 43.885 54.650 45.240 54.880 ;
        RECT 49.210 54.650 50.565 54.880 ;
        RECT 54.545 54.650 55.900 54.880 ;
        RECT 59.870 54.650 61.225 54.880 ;
        RECT 65.205 54.650 66.560 54.880 ;
        RECT 70.530 54.650 71.885 54.880 ;
        RECT 75.865 54.650 77.220 54.880 ;
        RECT 81.190 54.650 82.545 54.880 ;
        RECT 86.525 54.650 87.880 54.880 ;
        RECT 91.850 54.650 93.205 54.880 ;
        RECT 97.185 54.650 98.540 54.880 ;
        RECT 102.510 54.650 103.865 54.880 ;
        RECT 107.845 54.650 109.200 54.880 ;
        RECT 113.170 54.650 114.525 54.880 ;
        RECT 118.505 54.650 119.860 54.880 ;
        RECT 123.830 54.650 125.185 54.880 ;
        RECT 32.955 54.185 33.455 54.355 ;
        RECT 33.810 54.270 34.005 54.650 ;
        RECT 34.335 54.185 34.835 54.355 ;
        RECT 39.135 54.270 39.330 54.650 ;
        RECT 44.470 54.270 44.665 54.650 ;
        RECT 49.795 54.270 49.990 54.650 ;
        RECT 55.130 54.270 55.325 54.650 ;
        RECT 60.455 54.270 60.650 54.650 ;
        RECT 65.790 54.270 65.985 54.650 ;
        RECT 71.115 54.270 71.310 54.650 ;
        RECT 76.450 54.270 76.645 54.650 ;
        RECT 81.775 54.270 81.970 54.650 ;
        RECT 87.110 54.270 87.305 54.650 ;
        RECT 92.435 54.270 92.630 54.650 ;
        RECT 97.770 54.270 97.965 54.650 ;
        RECT 103.095 54.270 103.290 54.650 ;
        RECT 108.430 54.270 108.625 54.650 ;
        RECT 113.755 54.270 113.950 54.650 ;
        RECT 119.090 54.270 119.285 54.650 ;
        RECT 123.560 54.185 124.060 54.355 ;
        RECT 124.415 54.270 124.610 54.650 ;
        RECT 124.940 54.185 125.440 54.355 ;
        RECT 32.955 47.565 33.455 47.735 ;
        RECT 33.810 47.345 34.005 47.735 ;
        RECT 34.335 47.565 34.835 47.735 ;
        RECT 39.135 47.345 39.330 47.735 ;
        RECT 44.470 47.345 44.665 47.735 ;
        RECT 49.795 47.345 49.990 47.735 ;
        RECT 55.130 47.345 55.325 47.735 ;
        RECT 60.455 47.345 60.650 47.735 ;
        RECT 65.790 47.345 65.985 47.735 ;
        RECT 71.115 47.345 71.310 47.735 ;
        RECT 76.450 47.345 76.645 47.735 ;
        RECT 81.775 47.345 81.970 47.735 ;
        RECT 87.110 47.345 87.305 47.735 ;
        RECT 92.435 47.345 92.630 47.735 ;
        RECT 97.770 47.345 97.965 47.735 ;
        RECT 103.095 47.345 103.290 47.735 ;
        RECT 108.430 47.345 108.625 47.735 ;
        RECT 113.755 47.345 113.950 47.735 ;
        RECT 119.090 47.345 119.285 47.735 ;
        RECT 123.560 47.565 124.060 47.735 ;
        RECT 124.415 47.345 124.610 47.735 ;
        RECT 124.940 47.565 125.440 47.735 ;
        RECT 33.225 47.115 34.580 47.345 ;
        RECT 38.550 47.115 39.905 47.345 ;
        RECT 43.885 47.115 45.240 47.345 ;
        RECT 49.210 47.115 50.565 47.345 ;
        RECT 54.545 47.115 55.900 47.345 ;
        RECT 59.870 47.115 61.225 47.345 ;
        RECT 65.205 47.115 66.560 47.345 ;
        RECT 70.530 47.115 71.885 47.345 ;
        RECT 75.865 47.115 77.220 47.345 ;
        RECT 81.190 47.115 82.545 47.345 ;
        RECT 86.525 47.115 87.880 47.345 ;
        RECT 91.850 47.115 93.205 47.345 ;
        RECT 97.185 47.115 98.540 47.345 ;
        RECT 102.510 47.115 103.865 47.345 ;
        RECT 107.845 47.115 109.200 47.345 ;
        RECT 113.170 47.115 114.525 47.345 ;
        RECT 118.505 47.115 119.860 47.345 ;
        RECT 123.830 47.115 125.185 47.345 ;
        RECT 32.955 46.650 33.455 46.820 ;
        RECT 33.810 46.735 34.005 47.115 ;
        RECT 34.335 46.650 34.835 46.820 ;
        RECT 39.135 46.735 39.330 47.115 ;
        RECT 44.470 46.735 44.665 47.115 ;
        RECT 49.795 46.735 49.990 47.115 ;
        RECT 55.130 46.735 55.325 47.115 ;
        RECT 60.455 46.735 60.650 47.115 ;
        RECT 65.790 46.735 65.985 47.115 ;
        RECT 71.115 46.735 71.310 47.115 ;
        RECT 76.450 46.735 76.645 47.115 ;
        RECT 81.775 46.735 81.970 47.115 ;
        RECT 87.110 46.735 87.305 47.115 ;
        RECT 92.435 46.735 92.630 47.115 ;
        RECT 97.770 46.735 97.965 47.115 ;
        RECT 103.095 46.735 103.290 47.115 ;
        RECT 108.430 46.735 108.625 47.115 ;
        RECT 113.755 46.735 113.950 47.115 ;
        RECT 119.090 46.735 119.285 47.115 ;
        RECT 123.560 46.650 124.060 46.820 ;
        RECT 124.415 46.735 124.610 47.115 ;
        RECT 124.940 46.650 125.440 46.820 ;
        RECT 32.955 40.030 33.455 40.200 ;
        RECT 33.810 39.810 34.005 40.200 ;
        RECT 34.335 40.030 34.835 40.200 ;
        RECT 39.135 39.810 39.330 40.200 ;
        RECT 44.470 39.810 44.665 40.200 ;
        RECT 49.795 39.810 49.990 40.200 ;
        RECT 55.130 39.810 55.325 40.200 ;
        RECT 60.455 39.810 60.650 40.200 ;
        RECT 65.790 39.810 65.985 40.200 ;
        RECT 71.115 39.810 71.310 40.200 ;
        RECT 76.450 39.810 76.645 40.200 ;
        RECT 81.775 39.810 81.970 40.200 ;
        RECT 87.110 39.810 87.305 40.200 ;
        RECT 92.435 39.810 92.630 40.200 ;
        RECT 97.770 39.810 97.965 40.200 ;
        RECT 103.095 39.810 103.290 40.200 ;
        RECT 108.430 39.810 108.625 40.200 ;
        RECT 113.755 39.810 113.950 40.200 ;
        RECT 119.090 39.810 119.285 40.200 ;
        RECT 123.560 40.030 124.060 40.200 ;
        RECT 124.415 39.810 124.610 40.200 ;
        RECT 124.940 40.030 125.440 40.200 ;
        RECT 33.225 39.580 34.580 39.810 ;
        RECT 38.550 39.580 39.905 39.810 ;
        RECT 43.885 39.580 45.240 39.810 ;
        RECT 49.210 39.580 50.565 39.810 ;
        RECT 54.545 39.580 55.900 39.810 ;
        RECT 59.870 39.580 61.225 39.810 ;
        RECT 65.205 39.580 66.560 39.810 ;
        RECT 70.530 39.580 71.885 39.810 ;
        RECT 75.865 39.580 77.220 39.810 ;
        RECT 81.190 39.580 82.545 39.810 ;
        RECT 86.525 39.580 87.880 39.810 ;
        RECT 91.850 39.580 93.205 39.810 ;
        RECT 97.185 39.580 98.540 39.810 ;
        RECT 102.510 39.580 103.865 39.810 ;
        RECT 107.845 39.580 109.200 39.810 ;
        RECT 113.170 39.580 114.525 39.810 ;
        RECT 118.505 39.580 119.860 39.810 ;
        RECT 123.830 39.580 125.185 39.810 ;
        RECT 32.955 39.115 33.455 39.285 ;
        RECT 33.810 39.200 34.005 39.580 ;
        RECT 34.335 39.115 34.835 39.285 ;
        RECT 39.135 39.200 39.330 39.580 ;
        RECT 44.470 39.200 44.665 39.580 ;
        RECT 49.795 39.200 49.990 39.580 ;
        RECT 55.130 39.200 55.325 39.580 ;
        RECT 60.455 39.200 60.650 39.580 ;
        RECT 65.790 39.200 65.985 39.580 ;
        RECT 71.115 39.200 71.310 39.580 ;
        RECT 76.450 39.200 76.645 39.580 ;
        RECT 81.775 39.200 81.970 39.580 ;
        RECT 87.110 39.200 87.305 39.580 ;
        RECT 92.435 39.200 92.630 39.580 ;
        RECT 97.770 39.200 97.965 39.580 ;
        RECT 103.095 39.200 103.290 39.580 ;
        RECT 108.430 39.200 108.625 39.580 ;
        RECT 113.755 39.200 113.950 39.580 ;
        RECT 119.090 39.200 119.285 39.580 ;
        RECT 123.560 39.115 124.060 39.285 ;
        RECT 124.415 39.200 124.610 39.580 ;
        RECT 124.940 39.115 125.440 39.285 ;
        RECT 32.955 32.495 33.455 32.665 ;
        RECT 33.810 32.275 34.005 32.665 ;
        RECT 34.335 32.495 34.835 32.665 ;
        RECT 39.135 32.275 39.330 32.665 ;
        RECT 44.470 32.275 44.665 32.665 ;
        RECT 49.795 32.275 49.990 32.665 ;
        RECT 55.130 32.275 55.325 32.665 ;
        RECT 60.455 32.275 60.650 32.665 ;
        RECT 65.790 32.275 65.985 32.665 ;
        RECT 71.115 32.275 71.310 32.665 ;
        RECT 76.450 32.275 76.645 32.665 ;
        RECT 81.775 32.275 81.970 32.665 ;
        RECT 87.110 32.275 87.305 32.665 ;
        RECT 92.435 32.275 92.630 32.665 ;
        RECT 97.770 32.275 97.965 32.665 ;
        RECT 103.095 32.275 103.290 32.665 ;
        RECT 108.430 32.275 108.625 32.665 ;
        RECT 113.755 32.275 113.950 32.665 ;
        RECT 119.090 32.275 119.285 32.665 ;
        RECT 123.560 32.495 124.060 32.665 ;
        RECT 124.415 32.275 124.610 32.665 ;
        RECT 124.940 32.495 125.440 32.665 ;
        RECT 33.225 32.045 34.580 32.275 ;
        RECT 38.550 32.045 39.905 32.275 ;
        RECT 43.885 32.045 45.240 32.275 ;
        RECT 49.210 32.045 50.565 32.275 ;
        RECT 54.545 32.045 55.900 32.275 ;
        RECT 59.870 32.045 61.225 32.275 ;
        RECT 65.205 32.045 66.560 32.275 ;
        RECT 70.530 32.045 71.885 32.275 ;
        RECT 75.865 32.045 77.220 32.275 ;
        RECT 81.190 32.045 82.545 32.275 ;
        RECT 86.525 32.045 87.880 32.275 ;
        RECT 91.850 32.045 93.205 32.275 ;
        RECT 97.185 32.045 98.540 32.275 ;
        RECT 102.510 32.045 103.865 32.275 ;
        RECT 107.845 32.045 109.200 32.275 ;
        RECT 113.170 32.045 114.525 32.275 ;
        RECT 118.505 32.045 119.860 32.275 ;
        RECT 123.830 32.045 125.185 32.275 ;
        RECT 32.955 31.580 33.455 31.750 ;
        RECT 33.810 31.665 34.005 32.045 ;
        RECT 34.335 31.580 34.835 31.750 ;
        RECT 39.135 31.665 39.330 32.045 ;
        RECT 44.470 31.665 44.665 32.045 ;
        RECT 49.795 31.665 49.990 32.045 ;
        RECT 55.130 31.665 55.325 32.045 ;
        RECT 60.455 31.665 60.650 32.045 ;
        RECT 65.790 31.665 65.985 32.045 ;
        RECT 71.115 31.665 71.310 32.045 ;
        RECT 76.450 31.665 76.645 32.045 ;
        RECT 81.775 31.665 81.970 32.045 ;
        RECT 87.110 31.665 87.305 32.045 ;
        RECT 92.435 31.665 92.630 32.045 ;
        RECT 97.770 31.665 97.965 32.045 ;
        RECT 103.095 31.665 103.290 32.045 ;
        RECT 108.430 31.665 108.625 32.045 ;
        RECT 113.755 31.665 113.950 32.045 ;
        RECT 119.090 31.665 119.285 32.045 ;
        RECT 123.560 31.580 124.060 31.750 ;
        RECT 124.415 31.665 124.610 32.045 ;
        RECT 124.940 31.580 125.440 31.750 ;
        RECT 32.955 24.960 33.455 25.130 ;
        RECT 33.810 24.740 34.005 25.130 ;
        RECT 34.335 24.960 34.835 25.130 ;
        RECT 39.135 24.740 39.330 25.130 ;
        RECT 44.470 24.740 44.665 25.130 ;
        RECT 49.795 24.740 49.990 25.130 ;
        RECT 55.130 24.740 55.325 25.130 ;
        RECT 60.455 24.740 60.650 25.130 ;
        RECT 65.790 24.740 65.985 25.130 ;
        RECT 71.115 24.740 71.310 25.130 ;
        RECT 76.450 24.740 76.645 25.130 ;
        RECT 81.775 24.740 81.970 25.130 ;
        RECT 87.110 24.740 87.305 25.130 ;
        RECT 92.435 24.740 92.630 25.130 ;
        RECT 97.770 24.740 97.965 25.130 ;
        RECT 103.095 24.740 103.290 25.130 ;
        RECT 108.430 24.740 108.625 25.130 ;
        RECT 113.755 24.740 113.950 25.130 ;
        RECT 119.090 24.740 119.285 25.130 ;
        RECT 123.560 24.960 124.060 25.130 ;
        RECT 124.415 24.740 124.610 25.130 ;
        RECT 124.940 24.960 125.440 25.130 ;
        RECT 33.225 24.510 34.580 24.740 ;
        RECT 38.550 24.510 39.905 24.740 ;
        RECT 43.885 24.510 45.240 24.740 ;
        RECT 49.210 24.510 50.565 24.740 ;
        RECT 54.545 24.510 55.900 24.740 ;
        RECT 59.870 24.510 61.225 24.740 ;
        RECT 65.205 24.510 66.560 24.740 ;
        RECT 70.530 24.510 71.885 24.740 ;
        RECT 75.865 24.510 77.220 24.740 ;
        RECT 81.190 24.510 82.545 24.740 ;
        RECT 86.525 24.510 87.880 24.740 ;
        RECT 91.850 24.510 93.205 24.740 ;
        RECT 97.185 24.510 98.540 24.740 ;
        RECT 102.510 24.510 103.865 24.740 ;
        RECT 107.845 24.510 109.200 24.740 ;
        RECT 113.170 24.510 114.525 24.740 ;
        RECT 118.505 24.510 119.860 24.740 ;
        RECT 123.830 24.510 125.185 24.740 ;
        RECT 32.955 24.045 33.455 24.215 ;
        RECT 33.810 24.130 34.005 24.510 ;
        RECT 34.335 24.045 34.835 24.215 ;
        RECT 39.135 24.130 39.330 24.510 ;
        RECT 44.470 24.130 44.665 24.510 ;
        RECT 49.795 24.130 49.990 24.510 ;
        RECT 55.130 24.130 55.325 24.510 ;
        RECT 60.455 24.130 60.650 24.510 ;
        RECT 65.790 24.130 65.985 24.510 ;
        RECT 71.115 24.130 71.310 24.510 ;
        RECT 76.450 24.130 76.645 24.510 ;
        RECT 81.775 24.130 81.970 24.510 ;
        RECT 87.110 24.130 87.305 24.510 ;
        RECT 92.435 24.130 92.630 24.510 ;
        RECT 97.770 24.130 97.965 24.510 ;
        RECT 103.095 24.130 103.290 24.510 ;
        RECT 108.430 24.130 108.625 24.510 ;
        RECT 113.755 24.130 113.950 24.510 ;
        RECT 119.090 24.130 119.285 24.510 ;
        RECT 123.560 24.045 124.060 24.215 ;
        RECT 124.415 24.130 124.610 24.510 ;
        RECT 124.940 24.045 125.440 24.215 ;
        RECT 32.955 17.425 33.455 17.595 ;
        RECT 33.810 17.205 34.005 17.595 ;
        RECT 34.335 17.425 34.835 17.595 ;
        RECT 39.135 17.205 39.330 17.595 ;
        RECT 44.470 17.205 44.665 17.595 ;
        RECT 49.795 17.205 49.990 17.595 ;
        RECT 55.130 17.205 55.325 17.595 ;
        RECT 60.455 17.205 60.650 17.595 ;
        RECT 65.790 17.205 65.985 17.595 ;
        RECT 71.115 17.205 71.310 17.595 ;
        RECT 76.450 17.205 76.645 17.595 ;
        RECT 81.775 17.205 81.970 17.595 ;
        RECT 87.110 17.205 87.305 17.595 ;
        RECT 92.435 17.205 92.630 17.595 ;
        RECT 97.770 17.205 97.965 17.595 ;
        RECT 103.095 17.205 103.290 17.595 ;
        RECT 108.430 17.205 108.625 17.595 ;
        RECT 113.755 17.205 113.950 17.595 ;
        RECT 119.090 17.205 119.285 17.595 ;
        RECT 123.560 17.425 124.060 17.595 ;
        RECT 124.415 17.205 124.610 17.595 ;
        RECT 124.940 17.425 125.440 17.595 ;
        RECT 33.225 16.975 34.580 17.205 ;
        RECT 38.550 16.975 39.905 17.205 ;
        RECT 43.885 16.975 45.240 17.205 ;
        RECT 49.210 16.975 50.565 17.205 ;
        RECT 54.545 16.975 55.900 17.205 ;
        RECT 59.870 16.975 61.225 17.205 ;
        RECT 65.205 16.975 66.560 17.205 ;
        RECT 70.530 16.975 71.885 17.205 ;
        RECT 75.865 16.975 77.220 17.205 ;
        RECT 81.190 16.975 82.545 17.205 ;
        RECT 86.525 16.975 87.880 17.205 ;
        RECT 91.850 16.975 93.205 17.205 ;
        RECT 97.185 16.975 98.540 17.205 ;
        RECT 102.510 16.975 103.865 17.205 ;
        RECT 107.845 16.975 109.200 17.205 ;
        RECT 113.170 16.975 114.525 17.205 ;
        RECT 118.505 16.975 119.860 17.205 ;
        RECT 123.830 16.975 125.185 17.205 ;
        RECT 32.955 16.510 33.455 16.680 ;
        RECT 33.810 16.595 34.005 16.975 ;
        RECT 34.335 16.510 34.835 16.680 ;
        RECT 39.135 16.595 39.330 16.975 ;
        RECT 44.470 16.595 44.665 16.975 ;
        RECT 49.795 16.595 49.990 16.975 ;
        RECT 55.130 16.595 55.325 16.975 ;
        RECT 60.455 16.595 60.650 16.975 ;
        RECT 65.790 16.595 65.985 16.975 ;
        RECT 71.115 16.595 71.310 16.975 ;
        RECT 76.450 16.595 76.645 16.975 ;
        RECT 81.775 16.595 81.970 16.975 ;
        RECT 87.110 16.595 87.305 16.975 ;
        RECT 92.435 16.595 92.630 16.975 ;
        RECT 97.770 16.595 97.965 16.975 ;
        RECT 103.095 16.595 103.290 16.975 ;
        RECT 108.430 16.595 108.625 16.975 ;
        RECT 113.755 16.595 113.950 16.975 ;
        RECT 119.090 16.595 119.285 16.975 ;
        RECT 123.560 16.510 124.060 16.680 ;
        RECT 124.415 16.595 124.610 16.975 ;
        RECT 124.940 16.510 125.440 16.680 ;
        RECT 32.955 9.890 33.455 10.060 ;
        RECT 33.810 9.670 34.005 10.060 ;
        RECT 34.335 9.890 34.835 10.060 ;
        RECT 39.135 9.670 39.330 10.060 ;
        RECT 44.470 9.670 44.665 10.060 ;
        RECT 49.795 9.670 49.990 10.060 ;
        RECT 55.130 9.670 55.325 10.060 ;
        RECT 60.455 9.670 60.650 10.060 ;
        RECT 65.790 9.670 65.985 10.060 ;
        RECT 71.115 9.670 71.310 10.060 ;
        RECT 76.450 9.670 76.645 10.060 ;
        RECT 81.775 9.670 81.970 10.060 ;
        RECT 87.110 9.670 87.305 10.060 ;
        RECT 92.435 9.670 92.630 10.060 ;
        RECT 97.770 9.670 97.965 10.060 ;
        RECT 103.095 9.670 103.290 10.060 ;
        RECT 108.430 9.670 108.625 10.060 ;
        RECT 113.755 9.670 113.950 10.060 ;
        RECT 119.090 9.670 119.285 10.060 ;
        RECT 123.560 9.890 124.060 10.060 ;
        RECT 124.415 9.670 124.610 10.060 ;
        RECT 124.940 9.890 125.440 10.060 ;
        RECT 33.225 9.440 34.580 9.670 ;
        RECT 38.550 9.440 39.905 9.670 ;
        RECT 43.885 9.440 45.240 9.670 ;
        RECT 49.210 9.440 50.565 9.670 ;
        RECT 54.545 9.440 55.900 9.670 ;
        RECT 59.870 9.440 61.225 9.670 ;
        RECT 65.205 9.440 66.560 9.670 ;
        RECT 70.530 9.440 71.885 9.670 ;
        RECT 75.865 9.440 77.220 9.670 ;
        RECT 81.190 9.440 82.545 9.670 ;
        RECT 86.525 9.440 87.880 9.670 ;
        RECT 91.850 9.440 93.205 9.670 ;
        RECT 97.185 9.440 98.540 9.670 ;
        RECT 102.510 9.440 103.865 9.670 ;
        RECT 107.845 9.440 109.200 9.670 ;
        RECT 113.170 9.440 114.525 9.670 ;
        RECT 118.505 9.440 119.860 9.670 ;
        RECT 123.830 9.440 125.185 9.670 ;
        RECT 32.955 8.975 33.455 9.145 ;
        RECT 33.810 9.060 34.005 9.440 ;
        RECT 34.335 8.975 34.835 9.145 ;
        RECT 38.280 8.975 38.780 9.145 ;
        RECT 39.135 9.060 39.330 9.440 ;
        RECT 39.660 8.975 40.160 9.145 ;
        RECT 43.615 8.975 44.115 9.145 ;
        RECT 44.470 9.060 44.665 9.440 ;
        RECT 44.995 8.975 45.495 9.145 ;
        RECT 48.940 8.975 49.440 9.145 ;
        RECT 49.795 9.060 49.990 9.440 ;
        RECT 50.320 8.975 50.820 9.145 ;
        RECT 54.275 8.975 54.775 9.145 ;
        RECT 55.130 9.060 55.325 9.440 ;
        RECT 55.655 8.975 56.155 9.145 ;
        RECT 59.600 8.975 60.100 9.145 ;
        RECT 60.455 9.060 60.650 9.440 ;
        RECT 60.980 8.975 61.480 9.145 ;
        RECT 64.935 8.975 65.435 9.145 ;
        RECT 65.790 9.060 65.985 9.440 ;
        RECT 66.315 8.975 66.815 9.145 ;
        RECT 70.260 8.975 70.760 9.145 ;
        RECT 71.115 9.060 71.310 9.440 ;
        RECT 71.640 8.975 72.140 9.145 ;
        RECT 75.595 8.975 76.095 9.145 ;
        RECT 76.450 9.060 76.645 9.440 ;
        RECT 76.975 8.975 77.475 9.145 ;
        RECT 80.920 8.975 81.420 9.145 ;
        RECT 81.775 9.060 81.970 9.440 ;
        RECT 82.300 8.975 82.800 9.145 ;
        RECT 86.255 8.975 86.755 9.145 ;
        RECT 87.110 9.060 87.305 9.440 ;
        RECT 87.635 8.975 88.135 9.145 ;
        RECT 91.580 8.975 92.080 9.145 ;
        RECT 92.435 9.060 92.630 9.440 ;
        RECT 92.960 8.975 93.460 9.145 ;
        RECT 96.915 8.975 97.415 9.145 ;
        RECT 97.770 9.060 97.965 9.440 ;
        RECT 98.295 8.975 98.795 9.145 ;
        RECT 102.240 8.975 102.740 9.145 ;
        RECT 103.095 9.060 103.290 9.440 ;
        RECT 103.620 8.975 104.120 9.145 ;
        RECT 107.575 8.975 108.075 9.145 ;
        RECT 108.430 9.060 108.625 9.440 ;
        RECT 108.955 8.975 109.455 9.145 ;
        RECT 112.900 8.975 113.400 9.145 ;
        RECT 113.755 9.060 113.950 9.440 ;
        RECT 114.280 8.975 114.780 9.145 ;
        RECT 118.235 8.975 118.735 9.145 ;
        RECT 119.090 9.060 119.285 9.440 ;
        RECT 119.615 8.975 120.115 9.145 ;
        RECT 123.560 8.975 124.060 9.145 ;
        RECT 124.415 9.060 124.610 9.440 ;
        RECT 124.940 8.975 125.440 9.145 ;
        RECT 32.955 2.355 33.455 2.525 ;
        RECT 33.810 2.135 34.005 2.525 ;
        RECT 34.335 2.355 34.835 2.525 ;
        RECT 38.280 2.355 38.780 2.525 ;
        RECT 39.135 2.135 39.330 2.525 ;
        RECT 39.660 2.355 40.160 2.525 ;
        RECT 43.615 2.355 44.115 2.525 ;
        RECT 44.470 2.135 44.665 2.525 ;
        RECT 44.995 2.355 45.495 2.525 ;
        RECT 48.940 2.355 49.440 2.525 ;
        RECT 49.795 2.135 49.990 2.525 ;
        RECT 50.320 2.355 50.820 2.525 ;
        RECT 54.275 2.355 54.775 2.525 ;
        RECT 55.130 2.135 55.325 2.525 ;
        RECT 55.655 2.355 56.155 2.525 ;
        RECT 59.600 2.355 60.100 2.525 ;
        RECT 60.455 2.135 60.650 2.525 ;
        RECT 60.980 2.355 61.480 2.525 ;
        RECT 64.935 2.355 65.435 2.525 ;
        RECT 65.790 2.135 65.985 2.525 ;
        RECT 66.315 2.355 66.815 2.525 ;
        RECT 70.260 2.355 70.760 2.525 ;
        RECT 71.115 2.135 71.310 2.525 ;
        RECT 71.640 2.355 72.140 2.525 ;
        RECT 75.595 2.355 76.095 2.525 ;
        RECT 76.450 2.135 76.645 2.525 ;
        RECT 76.975 2.355 77.475 2.525 ;
        RECT 80.920 2.355 81.420 2.525 ;
        RECT 81.775 2.135 81.970 2.525 ;
        RECT 82.300 2.355 82.800 2.525 ;
        RECT 86.255 2.355 86.755 2.525 ;
        RECT 87.110 2.135 87.305 2.525 ;
        RECT 87.635 2.355 88.135 2.525 ;
        RECT 91.580 2.355 92.080 2.525 ;
        RECT 92.435 2.135 92.630 2.525 ;
        RECT 92.960 2.355 93.460 2.525 ;
        RECT 96.915 2.355 97.415 2.525 ;
        RECT 97.770 2.135 97.965 2.525 ;
        RECT 98.295 2.355 98.795 2.525 ;
        RECT 102.240 2.355 102.740 2.525 ;
        RECT 103.095 2.135 103.290 2.525 ;
        RECT 103.620 2.355 104.120 2.525 ;
        RECT 107.575 2.355 108.075 2.525 ;
        RECT 108.430 2.135 108.625 2.525 ;
        RECT 108.955 2.355 109.455 2.525 ;
        RECT 112.900 2.355 113.400 2.525 ;
        RECT 113.755 2.135 113.950 2.525 ;
        RECT 114.280 2.355 114.780 2.525 ;
        RECT 118.235 2.355 118.735 2.525 ;
        RECT 119.090 2.135 119.285 2.525 ;
        RECT 119.615 2.355 120.115 2.525 ;
        RECT 123.560 2.355 124.060 2.525 ;
        RECT 124.415 2.135 124.610 2.525 ;
        RECT 124.940 2.355 125.440 2.525 ;
        RECT 33.225 1.905 34.580 2.135 ;
        RECT 38.550 1.905 39.905 2.135 ;
        RECT 43.885 1.905 45.240 2.135 ;
        RECT 49.210 1.905 50.565 2.135 ;
        RECT 54.545 1.905 55.900 2.135 ;
        RECT 59.870 1.905 61.225 2.135 ;
        RECT 65.205 1.905 66.560 2.135 ;
        RECT 70.530 1.905 71.885 2.135 ;
        RECT 75.865 1.905 77.220 2.135 ;
        RECT 81.190 1.905 82.545 2.135 ;
        RECT 86.525 1.905 87.880 2.135 ;
        RECT 91.850 1.905 93.205 2.135 ;
        RECT 97.185 1.905 98.540 2.135 ;
        RECT 102.510 1.905 103.865 2.135 ;
        RECT 107.845 1.905 109.200 2.135 ;
        RECT 113.170 1.905 114.525 2.135 ;
        RECT 118.505 1.905 119.860 2.135 ;
        RECT 123.830 1.905 125.185 2.135 ;
        RECT 129.095 0.600 129.265 78.790 ;
        RECT 29.160 0.430 129.265 0.600 ;
      LAYER met1 ;
        RECT 29.060 78.690 129.365 79.060 ;
        RECT 0.330 62.175 21.930 63.425 ;
        RECT 0.330 54.035 21.930 55.285 ;
        RECT 0.330 45.895 21.930 47.145 ;
        RECT 0.330 37.755 21.930 39.005 ;
        RECT 0.330 29.615 21.930 30.865 ;
        RECT 0.330 21.475 21.930 22.725 ;
        RECT 0.330 13.335 21.930 14.585 ;
        RECT 0.330 5.195 21.930 6.445 ;
        RECT 29.060 0.700 29.430 78.690 ;
        RECT 128.995 78.255 129.365 78.690 ;
        RECT 32.195 76.760 33.435 76.990 ;
        RECT 33.745 76.810 34.070 77.375 ;
        RECT 34.355 76.760 35.545 76.990 ;
        RECT 32.195 76.335 32.455 76.760 ;
        RECT 35.285 75.685 35.545 76.760 ;
        RECT 37.520 76.760 38.760 76.990 ;
        RECT 39.070 76.810 39.395 77.375 ;
        RECT 39.680 76.760 40.870 76.990 ;
        RECT 37.520 76.335 37.780 76.760 ;
        RECT 40.610 75.685 40.870 76.760 ;
        RECT 42.855 76.760 44.095 76.990 ;
        RECT 44.405 76.810 44.730 77.375 ;
        RECT 45.015 76.760 46.205 76.990 ;
        RECT 42.855 76.335 43.115 76.760 ;
        RECT 45.945 75.685 46.205 76.760 ;
        RECT 48.180 76.760 49.420 76.990 ;
        RECT 49.730 76.810 50.055 77.375 ;
        RECT 50.340 76.760 51.530 76.990 ;
        RECT 48.180 76.335 48.440 76.760 ;
        RECT 51.270 75.685 51.530 76.760 ;
        RECT 53.515 76.760 54.755 76.990 ;
        RECT 55.065 76.810 55.390 77.375 ;
        RECT 55.675 76.760 56.865 76.990 ;
        RECT 53.515 76.335 53.775 76.760 ;
        RECT 56.605 75.685 56.865 76.760 ;
        RECT 58.840 76.760 60.080 76.990 ;
        RECT 60.390 76.810 60.715 77.375 ;
        RECT 61.000 76.760 62.190 76.990 ;
        RECT 58.840 76.335 59.100 76.760 ;
        RECT 61.930 75.685 62.190 76.760 ;
        RECT 64.175 76.760 65.415 76.990 ;
        RECT 65.725 76.810 66.050 77.375 ;
        RECT 66.335 76.760 67.525 76.990 ;
        RECT 64.175 76.335 64.435 76.760 ;
        RECT 67.265 75.685 67.525 76.760 ;
        RECT 69.500 76.760 70.740 76.990 ;
        RECT 71.050 76.810 71.375 77.375 ;
        RECT 71.660 76.760 72.850 76.990 ;
        RECT 69.500 76.335 69.760 76.760 ;
        RECT 72.590 75.685 72.850 76.760 ;
        RECT 74.835 76.760 76.075 76.990 ;
        RECT 76.385 76.810 76.710 77.375 ;
        RECT 76.995 76.760 78.185 76.990 ;
        RECT 74.835 76.335 75.095 76.760 ;
        RECT 77.925 75.685 78.185 76.760 ;
        RECT 80.160 76.760 81.400 76.990 ;
        RECT 81.710 76.810 82.035 77.375 ;
        RECT 82.320 76.760 83.510 76.990 ;
        RECT 80.160 76.335 80.420 76.760 ;
        RECT 83.250 75.685 83.510 76.760 ;
        RECT 85.495 76.760 86.735 76.990 ;
        RECT 87.045 76.810 87.370 77.375 ;
        RECT 87.655 76.760 88.845 76.990 ;
        RECT 85.495 76.335 85.755 76.760 ;
        RECT 88.585 75.685 88.845 76.760 ;
        RECT 90.820 76.760 92.060 76.990 ;
        RECT 92.370 76.810 92.695 77.375 ;
        RECT 92.980 76.760 94.170 76.990 ;
        RECT 90.820 76.335 91.080 76.760 ;
        RECT 93.910 75.685 94.170 76.760 ;
        RECT 96.155 76.760 97.395 76.990 ;
        RECT 97.705 76.810 98.030 77.375 ;
        RECT 98.315 76.760 99.505 76.990 ;
        RECT 96.155 76.335 96.415 76.760 ;
        RECT 99.245 75.685 99.505 76.760 ;
        RECT 101.480 76.760 102.720 76.990 ;
        RECT 103.030 76.810 103.355 77.375 ;
        RECT 103.640 76.760 104.830 76.990 ;
        RECT 101.480 76.335 101.740 76.760 ;
        RECT 104.570 75.685 104.830 76.760 ;
        RECT 106.815 76.760 108.055 76.990 ;
        RECT 108.365 76.810 108.690 77.375 ;
        RECT 108.975 76.760 110.165 76.990 ;
        RECT 106.815 76.335 107.075 76.760 ;
        RECT 109.905 75.685 110.165 76.760 ;
        RECT 112.140 76.760 113.380 76.990 ;
        RECT 113.690 76.810 114.015 77.375 ;
        RECT 114.300 76.760 115.490 76.990 ;
        RECT 112.140 76.335 112.400 76.760 ;
        RECT 115.230 75.685 115.490 76.760 ;
        RECT 117.475 76.760 118.715 76.990 ;
        RECT 119.025 76.810 119.350 77.375 ;
        RECT 119.635 76.760 120.825 76.990 ;
        RECT 117.475 76.335 117.735 76.760 ;
        RECT 120.565 75.685 120.825 76.760 ;
        RECT 122.800 76.760 124.040 76.990 ;
        RECT 124.350 76.810 124.675 77.375 ;
        RECT 124.960 76.760 126.150 76.990 ;
        RECT 122.800 76.335 123.060 76.760 ;
        RECT 125.890 75.685 126.150 76.760 ;
        RECT 32.245 70.370 32.505 71.505 ;
        RECT 32.245 70.140 33.435 70.370 ;
        RECT 32.195 69.225 33.435 69.455 ;
        RECT 33.745 69.275 34.070 70.405 ;
        RECT 35.335 70.370 35.595 70.875 ;
        RECT 34.355 70.140 35.595 70.370 ;
        RECT 37.570 70.370 37.830 71.505 ;
        RECT 37.570 70.140 38.760 70.370 ;
        RECT 34.355 69.225 35.545 69.455 ;
        RECT 39.070 69.275 39.395 70.405 ;
        RECT 40.660 70.370 40.920 70.875 ;
        RECT 39.680 70.140 40.920 70.370 ;
        RECT 42.905 70.370 43.165 71.505 ;
        RECT 42.905 70.140 44.095 70.370 ;
        RECT 44.405 69.275 44.730 70.405 ;
        RECT 45.995 70.370 46.255 70.875 ;
        RECT 45.015 70.140 46.255 70.370 ;
        RECT 48.230 70.370 48.490 71.505 ;
        RECT 48.230 70.140 49.420 70.370 ;
        RECT 49.730 69.275 50.055 70.405 ;
        RECT 51.320 70.370 51.580 70.875 ;
        RECT 50.340 70.140 51.580 70.370 ;
        RECT 53.565 70.370 53.825 71.505 ;
        RECT 53.565 70.140 54.755 70.370 ;
        RECT 55.065 69.275 55.390 70.405 ;
        RECT 56.655 70.370 56.915 70.875 ;
        RECT 55.675 70.140 56.915 70.370 ;
        RECT 58.890 70.370 59.150 71.505 ;
        RECT 58.890 70.140 60.080 70.370 ;
        RECT 60.390 69.275 60.715 70.405 ;
        RECT 61.980 70.370 62.240 70.875 ;
        RECT 61.000 70.140 62.240 70.370 ;
        RECT 64.225 70.370 64.485 71.505 ;
        RECT 64.225 70.140 65.415 70.370 ;
        RECT 65.725 69.275 66.050 70.405 ;
        RECT 67.315 70.370 67.575 70.875 ;
        RECT 66.335 70.140 67.575 70.370 ;
        RECT 69.550 70.370 69.810 71.505 ;
        RECT 69.550 70.140 70.740 70.370 ;
        RECT 71.050 69.275 71.375 70.405 ;
        RECT 72.640 70.370 72.900 70.875 ;
        RECT 71.660 70.140 72.900 70.370 ;
        RECT 74.885 70.370 75.145 71.505 ;
        RECT 74.885 70.140 76.075 70.370 ;
        RECT 32.195 68.800 32.455 69.225 ;
        RECT 35.285 68.150 35.545 69.225 ;
        RECT 74.835 69.225 76.075 69.455 ;
        RECT 76.385 69.275 76.710 70.405 ;
        RECT 77.975 70.370 78.235 70.875 ;
        RECT 76.995 70.140 78.235 70.370 ;
        RECT 80.210 70.370 80.470 71.505 ;
        RECT 80.210 70.140 81.400 70.370 ;
        RECT 81.710 69.275 82.035 70.405 ;
        RECT 83.300 70.370 83.560 70.875 ;
        RECT 82.320 70.140 83.560 70.370 ;
        RECT 85.545 70.370 85.805 71.505 ;
        RECT 85.545 70.140 86.735 70.370 ;
        RECT 87.045 69.275 87.370 70.405 ;
        RECT 88.635 70.370 88.895 70.875 ;
        RECT 87.655 70.140 88.895 70.370 ;
        RECT 90.870 70.370 91.130 71.505 ;
        RECT 90.870 70.140 92.060 70.370 ;
        RECT 92.370 69.275 92.695 70.405 ;
        RECT 93.960 70.370 94.220 70.875 ;
        RECT 92.980 70.140 94.220 70.370 ;
        RECT 96.205 70.370 96.465 71.505 ;
        RECT 96.205 70.140 97.395 70.370 ;
        RECT 97.705 69.275 98.030 70.405 ;
        RECT 99.295 70.370 99.555 70.875 ;
        RECT 98.315 70.140 99.555 70.370 ;
        RECT 101.530 70.370 101.790 71.505 ;
        RECT 101.530 70.140 102.720 70.370 ;
        RECT 103.030 69.275 103.355 70.405 ;
        RECT 104.620 70.370 104.880 70.875 ;
        RECT 103.640 70.140 104.880 70.370 ;
        RECT 106.865 70.370 107.125 71.505 ;
        RECT 106.865 70.140 108.055 70.370 ;
        RECT 108.365 69.275 108.690 70.405 ;
        RECT 109.955 70.370 110.215 70.875 ;
        RECT 108.975 70.140 110.215 70.370 ;
        RECT 112.190 70.370 112.450 71.505 ;
        RECT 112.190 70.140 113.380 70.370 ;
        RECT 113.690 69.275 114.015 70.405 ;
        RECT 115.280 70.370 115.540 70.875 ;
        RECT 114.300 70.140 115.540 70.370 ;
        RECT 117.525 70.370 117.785 71.505 ;
        RECT 117.525 70.140 118.715 70.370 ;
        RECT 117.475 69.225 118.715 69.455 ;
        RECT 119.025 69.275 119.350 70.405 ;
        RECT 120.615 70.370 120.875 70.875 ;
        RECT 119.635 70.140 120.875 70.370 ;
        RECT 122.850 70.370 123.110 71.505 ;
        RECT 122.850 70.140 124.040 70.370 ;
        RECT 122.800 69.225 124.040 69.455 ;
        RECT 124.350 69.275 124.675 70.405 ;
        RECT 125.940 70.370 126.200 70.875 ;
        RECT 124.960 70.140 126.200 70.370 ;
        RECT 124.960 69.225 126.150 69.455 ;
        RECT 74.835 68.800 75.095 69.225 ;
        RECT 117.475 68.800 117.735 69.225 ;
        RECT 122.800 68.800 123.060 69.225 ;
        RECT 125.890 68.150 126.150 69.225 ;
        RECT 32.245 62.835 32.505 63.970 ;
        RECT 32.245 62.605 33.435 62.835 ;
        RECT 32.195 61.690 33.435 61.920 ;
        RECT 33.745 61.740 34.070 62.870 ;
        RECT 35.335 62.835 35.595 63.340 ;
        RECT 34.355 62.605 35.595 62.835 ;
        RECT 34.355 61.690 35.545 61.920 ;
        RECT 39.070 61.740 39.395 62.870 ;
        RECT 44.405 61.740 44.730 62.870 ;
        RECT 49.730 61.740 50.055 62.870 ;
        RECT 55.065 61.740 55.390 62.870 ;
        RECT 60.390 61.740 60.715 62.870 ;
        RECT 65.725 61.740 66.050 62.870 ;
        RECT 71.050 61.740 71.375 62.870 ;
        RECT 76.385 61.740 76.710 62.870 ;
        RECT 81.710 61.740 82.035 62.870 ;
        RECT 87.045 61.740 87.370 62.870 ;
        RECT 92.370 61.740 92.695 62.870 ;
        RECT 97.705 61.740 98.030 62.870 ;
        RECT 103.030 61.740 103.355 62.870 ;
        RECT 108.365 61.740 108.690 62.870 ;
        RECT 113.690 61.740 114.015 62.870 ;
        RECT 119.025 61.740 119.350 62.870 ;
        RECT 122.850 62.835 123.110 63.970 ;
        RECT 122.850 62.605 124.040 62.835 ;
        RECT 32.195 61.265 32.455 61.690 ;
        RECT 35.285 60.615 35.545 61.690 ;
        RECT 122.800 61.690 124.040 61.920 ;
        RECT 124.350 61.740 124.675 62.870 ;
        RECT 125.940 62.835 126.200 63.340 ;
        RECT 124.960 62.605 126.200 62.835 ;
        RECT 124.960 61.690 126.150 61.920 ;
        RECT 122.800 61.265 123.060 61.690 ;
        RECT 125.890 60.615 126.150 61.690 ;
        RECT 32.245 55.300 32.505 56.435 ;
        RECT 32.245 55.070 33.435 55.300 ;
        RECT 32.195 54.155 33.435 54.385 ;
        RECT 33.745 54.205 34.070 55.335 ;
        RECT 35.335 55.300 35.595 55.805 ;
        RECT 34.355 55.070 35.595 55.300 ;
        RECT 34.355 54.155 35.545 54.385 ;
        RECT 39.070 54.205 39.395 55.335 ;
        RECT 44.405 54.205 44.730 55.335 ;
        RECT 49.730 54.205 50.055 55.335 ;
        RECT 55.065 54.205 55.390 55.335 ;
        RECT 60.390 54.205 60.715 55.335 ;
        RECT 65.725 54.205 66.050 55.335 ;
        RECT 71.050 54.205 71.375 55.335 ;
        RECT 76.385 54.205 76.710 55.335 ;
        RECT 81.710 54.205 82.035 55.335 ;
        RECT 87.045 54.205 87.370 55.335 ;
        RECT 92.370 54.205 92.695 55.335 ;
        RECT 97.705 54.205 98.030 55.335 ;
        RECT 103.030 54.205 103.355 55.335 ;
        RECT 108.365 54.205 108.690 55.335 ;
        RECT 113.690 54.205 114.015 55.335 ;
        RECT 119.025 54.205 119.350 55.335 ;
        RECT 122.850 55.300 123.110 56.435 ;
        RECT 122.850 55.070 124.040 55.300 ;
        RECT 32.195 53.730 32.455 54.155 ;
        RECT 35.285 53.080 35.545 54.155 ;
        RECT 122.800 54.155 124.040 54.385 ;
        RECT 124.350 54.205 124.675 55.335 ;
        RECT 125.940 55.300 126.200 55.805 ;
        RECT 124.960 55.070 126.200 55.300 ;
        RECT 124.960 54.155 126.150 54.385 ;
        RECT 122.800 53.730 123.060 54.155 ;
        RECT 125.890 53.080 126.150 54.155 ;
        RECT 32.245 47.765 32.505 48.900 ;
        RECT 32.245 47.535 33.435 47.765 ;
        RECT 32.195 46.620 33.435 46.850 ;
        RECT 33.745 46.670 34.070 47.800 ;
        RECT 35.335 47.765 35.595 48.270 ;
        RECT 34.355 47.535 35.595 47.765 ;
        RECT 34.355 46.620 35.545 46.850 ;
        RECT 39.070 46.670 39.395 47.800 ;
        RECT 44.405 46.670 44.730 47.800 ;
        RECT 49.730 46.670 50.055 47.800 ;
        RECT 55.065 46.670 55.390 47.800 ;
        RECT 60.390 46.670 60.715 47.800 ;
        RECT 65.725 46.670 66.050 47.800 ;
        RECT 71.050 46.670 71.375 47.800 ;
        RECT 76.385 46.670 76.710 47.800 ;
        RECT 81.710 46.670 82.035 47.800 ;
        RECT 87.045 46.670 87.370 47.800 ;
        RECT 92.370 46.670 92.695 47.800 ;
        RECT 97.705 46.670 98.030 47.800 ;
        RECT 103.030 46.670 103.355 47.800 ;
        RECT 108.365 46.670 108.690 47.800 ;
        RECT 113.690 46.670 114.015 47.800 ;
        RECT 119.025 46.670 119.350 47.800 ;
        RECT 122.850 47.765 123.110 48.900 ;
        RECT 122.850 47.535 124.040 47.765 ;
        RECT 32.195 46.195 32.455 46.620 ;
        RECT 35.285 45.545 35.545 46.620 ;
        RECT 122.800 46.620 124.040 46.850 ;
        RECT 124.350 46.670 124.675 47.800 ;
        RECT 125.940 47.765 126.200 48.270 ;
        RECT 124.960 47.535 126.200 47.765 ;
        RECT 124.960 46.620 126.150 46.850 ;
        RECT 122.800 46.195 123.060 46.620 ;
        RECT 125.890 45.545 126.150 46.620 ;
        RECT 32.245 40.230 32.505 41.365 ;
        RECT 32.245 40.000 33.435 40.230 ;
        RECT 32.195 39.085 33.435 39.315 ;
        RECT 33.745 39.135 34.070 40.265 ;
        RECT 35.335 40.230 35.595 40.735 ;
        RECT 34.355 40.000 35.595 40.230 ;
        RECT 34.355 39.085 35.545 39.315 ;
        RECT 39.070 39.135 39.395 40.265 ;
        RECT 44.405 39.135 44.730 40.265 ;
        RECT 49.730 39.135 50.055 40.265 ;
        RECT 55.065 39.135 55.390 40.265 ;
        RECT 60.390 39.135 60.715 40.265 ;
        RECT 65.725 39.135 66.050 40.265 ;
        RECT 71.050 39.135 71.375 40.265 ;
        RECT 76.385 39.135 76.710 40.265 ;
        RECT 81.710 39.135 82.035 40.265 ;
        RECT 87.045 39.135 87.370 40.265 ;
        RECT 92.370 39.135 92.695 40.265 ;
        RECT 97.705 39.135 98.030 40.265 ;
        RECT 103.030 39.135 103.355 40.265 ;
        RECT 108.365 39.135 108.690 40.265 ;
        RECT 113.690 39.135 114.015 40.265 ;
        RECT 119.025 39.135 119.350 40.265 ;
        RECT 122.850 40.230 123.110 41.365 ;
        RECT 122.850 40.000 124.040 40.230 ;
        RECT 32.195 38.660 32.455 39.085 ;
        RECT 35.285 38.010 35.545 39.085 ;
        RECT 122.800 39.085 124.040 39.315 ;
        RECT 124.350 39.135 124.675 40.265 ;
        RECT 125.940 40.230 126.200 40.735 ;
        RECT 124.960 40.000 126.200 40.230 ;
        RECT 124.960 39.085 126.150 39.315 ;
        RECT 122.800 38.660 123.060 39.085 ;
        RECT 125.890 38.010 126.150 39.085 ;
        RECT 32.245 32.695 32.505 33.830 ;
        RECT 32.245 32.465 33.435 32.695 ;
        RECT 32.195 31.550 33.435 31.780 ;
        RECT 33.745 31.600 34.070 32.730 ;
        RECT 35.335 32.695 35.595 33.200 ;
        RECT 34.355 32.465 35.595 32.695 ;
        RECT 34.355 31.550 35.545 31.780 ;
        RECT 39.070 31.600 39.395 32.730 ;
        RECT 44.405 31.600 44.730 32.730 ;
        RECT 49.730 31.600 50.055 32.730 ;
        RECT 55.065 31.600 55.390 32.730 ;
        RECT 60.390 31.600 60.715 32.730 ;
        RECT 65.725 31.600 66.050 32.730 ;
        RECT 71.050 31.600 71.375 32.730 ;
        RECT 76.385 31.600 76.710 32.730 ;
        RECT 81.710 31.600 82.035 32.730 ;
        RECT 87.045 31.600 87.370 32.730 ;
        RECT 92.370 31.600 92.695 32.730 ;
        RECT 97.705 31.600 98.030 32.730 ;
        RECT 103.030 31.600 103.355 32.730 ;
        RECT 108.365 31.600 108.690 32.730 ;
        RECT 113.690 31.600 114.015 32.730 ;
        RECT 119.025 31.600 119.350 32.730 ;
        RECT 122.850 32.695 123.110 33.830 ;
        RECT 122.850 32.465 124.040 32.695 ;
        RECT 32.195 31.125 32.455 31.550 ;
        RECT 35.285 30.475 35.545 31.550 ;
        RECT 122.800 31.550 124.040 31.780 ;
        RECT 124.350 31.600 124.675 32.730 ;
        RECT 125.940 32.695 126.200 33.200 ;
        RECT 124.960 32.465 126.200 32.695 ;
        RECT 124.960 31.550 126.150 31.780 ;
        RECT 122.800 31.125 123.060 31.550 ;
        RECT 125.890 30.475 126.150 31.550 ;
        RECT 32.245 25.160 32.505 26.295 ;
        RECT 32.245 24.930 33.435 25.160 ;
        RECT 32.195 24.015 33.435 24.245 ;
        RECT 33.745 24.065 34.070 25.195 ;
        RECT 35.335 25.160 35.595 25.665 ;
        RECT 34.355 24.930 35.595 25.160 ;
        RECT 34.355 24.015 35.545 24.245 ;
        RECT 39.070 24.065 39.395 25.195 ;
        RECT 44.405 24.065 44.730 25.195 ;
        RECT 49.730 24.065 50.055 25.195 ;
        RECT 55.065 24.065 55.390 25.195 ;
        RECT 60.390 24.065 60.715 25.195 ;
        RECT 65.725 24.065 66.050 25.195 ;
        RECT 71.050 24.065 71.375 25.195 ;
        RECT 76.385 24.065 76.710 25.195 ;
        RECT 81.710 24.065 82.035 25.195 ;
        RECT 87.045 24.065 87.370 25.195 ;
        RECT 92.370 24.065 92.695 25.195 ;
        RECT 97.705 24.065 98.030 25.195 ;
        RECT 103.030 24.065 103.355 25.195 ;
        RECT 108.365 24.065 108.690 25.195 ;
        RECT 113.690 24.065 114.015 25.195 ;
        RECT 119.025 24.065 119.350 25.195 ;
        RECT 122.850 25.160 123.110 26.295 ;
        RECT 122.850 24.930 124.040 25.160 ;
        RECT 32.195 23.590 32.455 24.015 ;
        RECT 35.285 22.940 35.545 24.015 ;
        RECT 122.800 24.015 124.040 24.245 ;
        RECT 124.350 24.065 124.675 25.195 ;
        RECT 125.940 25.160 126.200 25.665 ;
        RECT 124.960 24.930 126.200 25.160 ;
        RECT 124.960 24.015 126.150 24.245 ;
        RECT 122.800 23.590 123.060 24.015 ;
        RECT 125.890 22.940 126.150 24.015 ;
        RECT 32.245 17.625 32.505 18.760 ;
        RECT 32.245 17.395 33.435 17.625 ;
        RECT 32.195 16.480 33.435 16.710 ;
        RECT 33.745 16.530 34.070 17.660 ;
        RECT 35.335 17.625 35.595 18.130 ;
        RECT 34.355 17.395 35.595 17.625 ;
        RECT 34.355 16.480 35.545 16.710 ;
        RECT 39.070 16.530 39.395 17.660 ;
        RECT 44.405 16.530 44.730 17.660 ;
        RECT 49.730 16.530 50.055 17.660 ;
        RECT 55.065 16.530 55.390 17.660 ;
        RECT 60.390 16.530 60.715 17.660 ;
        RECT 65.725 16.530 66.050 17.660 ;
        RECT 71.050 16.530 71.375 17.660 ;
        RECT 76.385 16.530 76.710 17.660 ;
        RECT 81.710 16.530 82.035 17.660 ;
        RECT 87.045 16.530 87.370 17.660 ;
        RECT 92.370 16.530 92.695 17.660 ;
        RECT 97.705 16.530 98.030 17.660 ;
        RECT 103.030 16.530 103.355 17.660 ;
        RECT 108.365 16.530 108.690 17.660 ;
        RECT 113.690 16.530 114.015 17.660 ;
        RECT 119.025 16.530 119.350 17.660 ;
        RECT 122.850 17.625 123.110 18.760 ;
        RECT 122.850 17.395 124.040 17.625 ;
        RECT 32.195 16.055 32.455 16.480 ;
        RECT 35.285 15.405 35.545 16.480 ;
        RECT 122.800 16.480 124.040 16.710 ;
        RECT 124.350 16.530 124.675 17.660 ;
        RECT 125.940 17.625 126.200 18.130 ;
        RECT 124.960 17.395 126.200 17.625 ;
        RECT 124.960 16.480 126.150 16.710 ;
        RECT 122.800 16.055 123.060 16.480 ;
        RECT 125.890 15.405 126.150 16.480 ;
        RECT 32.245 10.090 32.505 11.225 ;
        RECT 32.245 9.860 33.435 10.090 ;
        RECT 32.195 8.945 33.435 9.175 ;
        RECT 33.745 8.995 34.070 10.125 ;
        RECT 35.335 10.090 35.595 10.595 ;
        RECT 34.355 9.860 35.595 10.090 ;
        RECT 34.355 8.945 35.545 9.175 ;
        RECT 32.195 8.520 32.455 8.945 ;
        RECT 35.285 7.870 35.545 8.945 ;
        RECT 37.520 8.945 38.760 9.175 ;
        RECT 39.070 8.995 39.395 10.125 ;
        RECT 39.680 8.945 40.870 9.175 ;
        RECT 37.520 8.520 37.780 8.945 ;
        RECT 40.610 7.870 40.870 8.945 ;
        RECT 42.855 8.945 44.095 9.175 ;
        RECT 44.405 8.995 44.730 10.125 ;
        RECT 45.015 8.945 46.205 9.175 ;
        RECT 42.855 8.520 43.115 8.945 ;
        RECT 45.945 7.870 46.205 8.945 ;
        RECT 48.180 8.945 49.420 9.175 ;
        RECT 49.730 8.995 50.055 10.125 ;
        RECT 50.340 8.945 51.530 9.175 ;
        RECT 48.180 8.520 48.440 8.945 ;
        RECT 51.270 7.870 51.530 8.945 ;
        RECT 53.515 8.945 54.755 9.175 ;
        RECT 55.065 8.995 55.390 10.125 ;
        RECT 55.675 8.945 56.865 9.175 ;
        RECT 53.515 8.520 53.775 8.945 ;
        RECT 56.605 7.870 56.865 8.945 ;
        RECT 58.840 8.945 60.080 9.175 ;
        RECT 60.390 8.995 60.715 10.125 ;
        RECT 61.000 8.945 62.190 9.175 ;
        RECT 58.840 8.520 59.100 8.945 ;
        RECT 61.930 7.870 62.190 8.945 ;
        RECT 64.175 8.945 65.415 9.175 ;
        RECT 65.725 8.995 66.050 10.125 ;
        RECT 66.335 8.945 67.525 9.175 ;
        RECT 64.175 8.520 64.435 8.945 ;
        RECT 67.265 7.870 67.525 8.945 ;
        RECT 69.500 8.945 70.740 9.175 ;
        RECT 71.050 8.995 71.375 10.125 ;
        RECT 71.660 8.945 72.850 9.175 ;
        RECT 69.500 8.520 69.760 8.945 ;
        RECT 72.590 7.870 72.850 8.945 ;
        RECT 74.835 8.945 76.075 9.175 ;
        RECT 76.385 8.995 76.710 10.125 ;
        RECT 76.995 8.945 78.185 9.175 ;
        RECT 74.835 8.520 75.095 8.945 ;
        RECT 77.925 7.870 78.185 8.945 ;
        RECT 80.160 8.945 81.400 9.175 ;
        RECT 81.710 8.995 82.035 10.125 ;
        RECT 82.320 8.945 83.510 9.175 ;
        RECT 80.160 8.520 80.420 8.945 ;
        RECT 83.250 7.870 83.510 8.945 ;
        RECT 85.495 8.945 86.735 9.175 ;
        RECT 87.045 8.995 87.370 10.125 ;
        RECT 87.655 8.945 88.845 9.175 ;
        RECT 85.495 8.520 85.755 8.945 ;
        RECT 88.585 7.870 88.845 8.945 ;
        RECT 90.820 8.945 92.060 9.175 ;
        RECT 92.370 8.995 92.695 10.125 ;
        RECT 92.980 8.945 94.170 9.175 ;
        RECT 90.820 8.520 91.080 8.945 ;
        RECT 93.910 7.870 94.170 8.945 ;
        RECT 96.155 8.945 97.395 9.175 ;
        RECT 97.705 8.995 98.030 10.125 ;
        RECT 98.315 8.945 99.505 9.175 ;
        RECT 96.155 8.520 96.415 8.945 ;
        RECT 99.245 7.870 99.505 8.945 ;
        RECT 101.480 8.945 102.720 9.175 ;
        RECT 103.030 8.995 103.355 10.125 ;
        RECT 103.640 8.945 104.830 9.175 ;
        RECT 101.480 8.520 101.740 8.945 ;
        RECT 104.570 7.870 104.830 8.945 ;
        RECT 106.815 8.945 108.055 9.175 ;
        RECT 108.365 8.995 108.690 10.125 ;
        RECT 108.975 8.945 110.165 9.175 ;
        RECT 106.815 8.520 107.075 8.945 ;
        RECT 109.905 7.870 110.165 8.945 ;
        RECT 112.140 8.945 113.380 9.175 ;
        RECT 113.690 8.995 114.015 10.125 ;
        RECT 114.300 8.945 115.490 9.175 ;
        RECT 112.140 8.520 112.400 8.945 ;
        RECT 115.230 7.870 115.490 8.945 ;
        RECT 117.475 8.945 118.715 9.175 ;
        RECT 119.025 8.995 119.350 10.125 ;
        RECT 122.850 10.090 123.110 11.225 ;
        RECT 122.850 9.860 124.040 10.090 ;
        RECT 119.635 8.945 120.825 9.175 ;
        RECT 117.475 8.520 117.735 8.945 ;
        RECT 120.565 7.870 120.825 8.945 ;
        RECT 122.800 8.945 124.040 9.175 ;
        RECT 124.350 8.995 124.675 10.125 ;
        RECT 125.940 10.090 126.200 10.595 ;
        RECT 124.960 9.860 126.200 10.090 ;
        RECT 124.960 8.945 126.150 9.175 ;
        RECT 122.800 8.520 123.060 8.945 ;
        RECT 125.890 7.870 126.150 8.945 ;
        RECT 32.245 2.555 32.505 3.690 ;
        RECT 32.245 2.325 33.435 2.555 ;
        RECT 33.745 2.025 34.070 2.590 ;
        RECT 35.335 2.555 35.595 3.060 ;
        RECT 34.355 2.325 35.595 2.555 ;
        RECT 37.570 2.555 37.830 3.690 ;
        RECT 37.570 2.325 38.760 2.555 ;
        RECT 39.070 2.025 39.395 2.590 ;
        RECT 40.660 2.555 40.920 3.060 ;
        RECT 39.680 2.325 40.920 2.555 ;
        RECT 42.905 2.555 43.165 3.690 ;
        RECT 42.905 2.325 44.095 2.555 ;
        RECT 44.405 2.025 44.730 2.590 ;
        RECT 45.995 2.555 46.255 3.060 ;
        RECT 45.015 2.325 46.255 2.555 ;
        RECT 48.230 2.555 48.490 3.690 ;
        RECT 48.230 2.325 49.420 2.555 ;
        RECT 49.730 2.025 50.055 2.590 ;
        RECT 51.320 2.555 51.580 3.060 ;
        RECT 50.340 2.325 51.580 2.555 ;
        RECT 53.565 2.555 53.825 3.690 ;
        RECT 53.565 2.325 54.755 2.555 ;
        RECT 55.065 2.025 55.390 2.590 ;
        RECT 56.655 2.555 56.915 3.060 ;
        RECT 55.675 2.325 56.915 2.555 ;
        RECT 58.890 2.555 59.150 3.690 ;
        RECT 58.890 2.325 60.080 2.555 ;
        RECT 60.390 2.025 60.715 2.590 ;
        RECT 61.980 2.555 62.240 3.060 ;
        RECT 61.000 2.325 62.240 2.555 ;
        RECT 64.225 2.555 64.485 3.690 ;
        RECT 64.225 2.325 65.415 2.555 ;
        RECT 65.725 2.025 66.050 2.590 ;
        RECT 67.315 2.555 67.575 3.060 ;
        RECT 66.335 2.325 67.575 2.555 ;
        RECT 69.550 2.555 69.810 3.690 ;
        RECT 69.550 2.325 70.740 2.555 ;
        RECT 71.050 2.025 71.375 2.590 ;
        RECT 72.640 2.555 72.900 3.060 ;
        RECT 71.660 2.325 72.900 2.555 ;
        RECT 74.885 2.555 75.145 3.690 ;
        RECT 74.885 2.325 76.075 2.555 ;
        RECT 76.385 2.025 76.710 2.590 ;
        RECT 77.975 2.555 78.235 3.060 ;
        RECT 76.995 2.325 78.235 2.555 ;
        RECT 80.210 2.555 80.470 3.690 ;
        RECT 80.210 2.325 81.400 2.555 ;
        RECT 81.710 2.025 82.035 2.590 ;
        RECT 83.300 2.555 83.560 3.060 ;
        RECT 82.320 2.325 83.560 2.555 ;
        RECT 85.545 2.555 85.805 3.690 ;
        RECT 85.545 2.325 86.735 2.555 ;
        RECT 87.045 2.025 87.370 2.590 ;
        RECT 88.635 2.555 88.895 3.060 ;
        RECT 87.655 2.325 88.895 2.555 ;
        RECT 90.870 2.555 91.130 3.690 ;
        RECT 90.870 2.325 92.060 2.555 ;
        RECT 92.370 2.025 92.695 2.590 ;
        RECT 93.960 2.555 94.220 3.060 ;
        RECT 92.980 2.325 94.220 2.555 ;
        RECT 96.205 2.555 96.465 3.690 ;
        RECT 96.205 2.325 97.395 2.555 ;
        RECT 97.705 2.025 98.030 2.590 ;
        RECT 99.295 2.555 99.555 3.060 ;
        RECT 98.315 2.325 99.555 2.555 ;
        RECT 101.530 2.555 101.790 3.690 ;
        RECT 101.530 2.325 102.720 2.555 ;
        RECT 103.030 2.025 103.355 2.590 ;
        RECT 104.620 2.555 104.880 3.060 ;
        RECT 103.640 2.325 104.880 2.555 ;
        RECT 106.865 2.555 107.125 3.690 ;
        RECT 106.865 2.325 108.055 2.555 ;
        RECT 108.365 2.025 108.690 2.590 ;
        RECT 109.955 2.555 110.215 3.060 ;
        RECT 108.975 2.325 110.215 2.555 ;
        RECT 112.190 2.555 112.450 3.690 ;
        RECT 112.190 2.325 113.380 2.555 ;
        RECT 113.690 2.025 114.015 2.590 ;
        RECT 115.280 2.555 115.540 3.060 ;
        RECT 114.300 2.325 115.540 2.555 ;
        RECT 117.525 2.555 117.785 3.690 ;
        RECT 117.525 2.325 118.715 2.555 ;
        RECT 119.025 2.025 119.350 2.590 ;
        RECT 120.615 2.555 120.875 3.060 ;
        RECT 119.635 2.325 120.875 2.555 ;
        RECT 122.850 2.555 123.110 3.690 ;
        RECT 122.850 2.325 124.040 2.555 ;
        RECT 124.350 2.025 124.675 2.590 ;
        RECT 125.940 2.555 126.200 3.060 ;
        RECT 124.960 2.325 126.200 2.555 ;
        RECT 127.520 1.045 129.365 78.255 ;
        RECT 128.640 1.025 129.365 1.045 ;
        RECT 128.995 0.700 129.365 1.025 ;
        RECT 29.060 0.330 129.365 0.700 ;
      LAYER met2 ;
        RECT 78.955 81.440 107.070 84.510 ;
        RECT 74.790 81.430 107.070 81.440 ;
        RECT 74.755 81.150 107.070 81.430 ;
        RECT 125.740 81.310 128.670 84.505 ;
        RECT 74.790 81.140 107.070 81.150 ;
        RECT 127.520 78.255 128.660 81.310 ;
        RECT 31.240 76.815 128.660 78.255 ;
        RECT 31.465 76.645 31.835 76.655 ;
        RECT 32.195 76.645 32.455 76.815 ;
        RECT 31.465 76.385 32.485 76.645 ;
        RECT 31.465 76.375 31.835 76.385 ;
        RECT 35.285 75.995 35.545 76.815 ;
        RECT 36.790 76.645 37.160 76.655 ;
        RECT 37.520 76.645 37.780 76.815 ;
        RECT 36.790 76.385 37.810 76.645 ;
        RECT 36.790 76.375 37.160 76.385 ;
        RECT 35.960 75.995 36.330 76.005 ;
        RECT 40.610 75.995 40.870 76.815 ;
        RECT 42.125 76.645 42.495 76.655 ;
        RECT 42.855 76.645 43.115 76.815 ;
        RECT 42.125 76.385 43.145 76.645 ;
        RECT 42.125 76.375 42.495 76.385 ;
        RECT 41.285 75.995 41.655 76.005 ;
        RECT 45.945 75.995 46.205 76.815 ;
        RECT 47.450 76.645 47.820 76.655 ;
        RECT 48.180 76.645 48.440 76.815 ;
        RECT 47.450 76.385 48.470 76.645 ;
        RECT 47.450 76.375 47.820 76.385 ;
        RECT 46.620 75.995 46.990 76.005 ;
        RECT 51.270 75.995 51.530 76.815 ;
        RECT 52.785 76.645 53.155 76.655 ;
        RECT 53.515 76.645 53.775 76.815 ;
        RECT 52.785 76.385 53.805 76.645 ;
        RECT 52.785 76.375 53.155 76.385 ;
        RECT 51.945 75.995 52.315 76.005 ;
        RECT 56.605 75.995 56.865 76.815 ;
        RECT 58.110 76.645 58.480 76.655 ;
        RECT 58.840 76.645 59.100 76.815 ;
        RECT 58.110 76.385 59.130 76.645 ;
        RECT 58.110 76.375 58.480 76.385 ;
        RECT 57.280 75.995 57.650 76.005 ;
        RECT 61.930 75.995 62.190 76.815 ;
        RECT 63.445 76.645 63.815 76.655 ;
        RECT 64.175 76.645 64.435 76.815 ;
        RECT 63.445 76.385 64.465 76.645 ;
        RECT 63.445 76.375 63.815 76.385 ;
        RECT 62.605 75.995 62.975 76.005 ;
        RECT 67.265 75.995 67.525 76.815 ;
        RECT 68.770 76.645 69.140 76.655 ;
        RECT 69.500 76.645 69.760 76.815 ;
        RECT 68.770 76.385 69.790 76.645 ;
        RECT 68.770 76.375 69.140 76.385 ;
        RECT 67.940 75.995 68.310 76.005 ;
        RECT 72.590 75.995 72.850 76.815 ;
        RECT 74.105 76.645 74.475 76.655 ;
        RECT 74.835 76.645 75.095 76.815 ;
        RECT 74.105 76.385 75.125 76.645 ;
        RECT 74.105 76.375 74.475 76.385 ;
        RECT 73.265 75.995 73.635 76.005 ;
        RECT 77.925 75.995 78.185 76.815 ;
        RECT 79.430 76.645 79.800 76.655 ;
        RECT 80.160 76.645 80.420 76.815 ;
        RECT 79.430 76.385 80.450 76.645 ;
        RECT 79.430 76.375 79.800 76.385 ;
        RECT 78.600 75.995 78.970 76.005 ;
        RECT 83.250 75.995 83.510 76.815 ;
        RECT 84.765 76.645 85.135 76.655 ;
        RECT 85.495 76.645 85.755 76.815 ;
        RECT 84.765 76.385 85.785 76.645 ;
        RECT 84.765 76.375 85.135 76.385 ;
        RECT 83.925 75.995 84.295 76.005 ;
        RECT 88.585 75.995 88.845 76.815 ;
        RECT 90.090 76.645 90.460 76.655 ;
        RECT 90.820 76.645 91.080 76.815 ;
        RECT 90.090 76.385 91.110 76.645 ;
        RECT 90.090 76.375 90.460 76.385 ;
        RECT 89.260 75.995 89.630 76.005 ;
        RECT 93.910 75.995 94.170 76.815 ;
        RECT 95.425 76.645 95.795 76.655 ;
        RECT 96.155 76.645 96.415 76.815 ;
        RECT 95.425 76.385 96.445 76.645 ;
        RECT 95.425 76.375 95.795 76.385 ;
        RECT 94.585 75.995 94.955 76.005 ;
        RECT 99.245 75.995 99.505 76.815 ;
        RECT 100.750 76.645 101.120 76.655 ;
        RECT 101.480 76.645 101.740 76.815 ;
        RECT 100.750 76.385 101.770 76.645 ;
        RECT 100.750 76.375 101.120 76.385 ;
        RECT 99.920 75.995 100.290 76.005 ;
        RECT 104.570 75.995 104.830 76.815 ;
        RECT 106.085 76.645 106.455 76.655 ;
        RECT 106.815 76.645 107.075 76.815 ;
        RECT 106.085 76.385 107.105 76.645 ;
        RECT 106.085 76.375 106.455 76.385 ;
        RECT 105.245 75.995 105.615 76.005 ;
        RECT 109.905 75.995 110.165 76.815 ;
        RECT 111.410 76.645 111.780 76.655 ;
        RECT 112.140 76.645 112.400 76.815 ;
        RECT 111.410 76.385 112.430 76.645 ;
        RECT 111.410 76.375 111.780 76.385 ;
        RECT 110.580 75.995 110.950 76.005 ;
        RECT 115.230 75.995 115.490 76.815 ;
        RECT 116.745 76.645 117.115 76.655 ;
        RECT 117.475 76.645 117.735 76.815 ;
        RECT 116.745 76.385 117.765 76.645 ;
        RECT 116.745 76.375 117.115 76.385 ;
        RECT 115.905 75.995 116.275 76.005 ;
        RECT 120.565 75.995 120.825 76.815 ;
        RECT 122.070 76.645 122.440 76.655 ;
        RECT 122.800 76.645 123.060 76.815 ;
        RECT 122.070 76.385 123.090 76.645 ;
        RECT 122.070 76.375 122.440 76.385 ;
        RECT 121.240 75.995 121.610 76.005 ;
        RECT 125.890 75.995 126.150 76.815 ;
        RECT 126.565 75.995 126.935 76.005 ;
        RECT 35.255 75.735 36.330 75.995 ;
        RECT 40.580 75.735 41.655 75.995 ;
        RECT 45.915 75.735 46.990 75.995 ;
        RECT 51.240 75.735 52.315 75.995 ;
        RECT 56.575 75.735 57.650 75.995 ;
        RECT 61.900 75.735 62.975 75.995 ;
        RECT 67.235 75.735 68.310 75.995 ;
        RECT 72.560 75.735 73.635 75.995 ;
        RECT 77.895 75.735 78.970 75.995 ;
        RECT 83.220 75.735 84.295 75.995 ;
        RECT 88.555 75.735 89.630 75.995 ;
        RECT 93.880 75.735 94.955 75.995 ;
        RECT 99.215 75.735 100.290 75.995 ;
        RECT 104.540 75.735 105.615 75.995 ;
        RECT 109.875 75.735 110.950 75.995 ;
        RECT 115.200 75.735 116.275 75.995 ;
        RECT 120.535 75.735 121.610 75.995 ;
        RECT 125.860 75.735 126.935 75.995 ;
        RECT 35.960 75.725 36.330 75.735 ;
        RECT 41.285 75.725 41.655 75.735 ;
        RECT 46.620 75.725 46.990 75.735 ;
        RECT 51.945 75.725 52.315 75.735 ;
        RECT 57.280 75.725 57.650 75.735 ;
        RECT 62.605 75.725 62.975 75.735 ;
        RECT 67.940 75.725 68.310 75.735 ;
        RECT 73.265 75.725 73.635 75.735 ;
        RECT 78.600 75.725 78.970 75.735 ;
        RECT 83.925 75.725 84.295 75.735 ;
        RECT 89.260 75.725 89.630 75.735 ;
        RECT 94.585 75.725 94.955 75.735 ;
        RECT 99.920 75.725 100.290 75.735 ;
        RECT 105.245 75.725 105.615 75.735 ;
        RECT 110.580 75.725 110.950 75.735 ;
        RECT 115.905 75.725 116.275 75.735 ;
        RECT 121.240 75.725 121.610 75.735 ;
        RECT 126.565 75.725 126.935 75.735 ;
        RECT 4.215 1.535 6.110 71.635 ;
        RECT 18.215 1.535 20.110 71.635 ;
        RECT 31.460 71.475 31.830 71.485 ;
        RECT 36.785 71.475 37.155 71.485 ;
        RECT 42.120 71.475 42.490 71.485 ;
        RECT 47.445 71.475 47.815 71.485 ;
        RECT 52.780 71.475 53.150 71.485 ;
        RECT 58.105 71.475 58.475 71.485 ;
        RECT 63.440 71.475 63.810 71.485 ;
        RECT 68.765 71.475 69.135 71.485 ;
        RECT 74.100 71.475 74.470 71.485 ;
        RECT 79.425 71.475 79.795 71.485 ;
        RECT 84.760 71.475 85.130 71.485 ;
        RECT 90.085 71.475 90.455 71.485 ;
        RECT 95.420 71.475 95.790 71.485 ;
        RECT 100.745 71.475 101.115 71.485 ;
        RECT 106.080 71.475 106.450 71.485 ;
        RECT 111.405 71.475 111.775 71.485 ;
        RECT 116.740 71.475 117.110 71.485 ;
        RECT 122.065 71.475 122.435 71.485 ;
        RECT 31.460 71.215 32.535 71.475 ;
        RECT 36.785 71.215 37.860 71.475 ;
        RECT 42.120 71.215 43.195 71.475 ;
        RECT 47.445 71.215 48.520 71.475 ;
        RECT 52.780 71.215 53.855 71.475 ;
        RECT 58.105 71.215 59.180 71.475 ;
        RECT 63.440 71.215 64.515 71.475 ;
        RECT 68.765 71.215 69.840 71.475 ;
        RECT 74.100 71.215 75.175 71.475 ;
        RECT 79.425 71.215 80.500 71.475 ;
        RECT 84.760 71.215 85.835 71.475 ;
        RECT 90.085 71.215 91.160 71.475 ;
        RECT 95.420 71.215 96.495 71.475 ;
        RECT 100.745 71.215 101.820 71.475 ;
        RECT 106.080 71.215 107.155 71.475 ;
        RECT 111.405 71.215 112.480 71.475 ;
        RECT 116.740 71.215 117.815 71.475 ;
        RECT 122.065 71.215 123.140 71.475 ;
        RECT 31.460 71.205 31.830 71.215 ;
        RECT 32.245 70.405 32.505 71.215 ;
        RECT 36.785 71.205 37.155 71.215 ;
        RECT 35.965 70.845 36.335 70.855 ;
        RECT 35.305 70.585 36.335 70.845 ;
        RECT 35.335 70.405 35.595 70.585 ;
        RECT 35.965 70.575 36.335 70.585 ;
        RECT 37.570 70.405 37.830 71.215 ;
        RECT 42.120 71.205 42.490 71.215 ;
        RECT 41.290 70.845 41.660 70.855 ;
        RECT 40.630 70.585 41.660 70.845 ;
        RECT 40.660 70.405 40.920 70.585 ;
        RECT 41.290 70.575 41.660 70.585 ;
        RECT 42.905 70.405 43.165 71.215 ;
        RECT 47.445 71.205 47.815 71.215 ;
        RECT 46.625 70.845 46.995 70.855 ;
        RECT 45.965 70.585 46.995 70.845 ;
        RECT 45.995 70.405 46.255 70.585 ;
        RECT 46.625 70.575 46.995 70.585 ;
        RECT 48.230 70.405 48.490 71.215 ;
        RECT 52.780 71.205 53.150 71.215 ;
        RECT 51.950 70.845 52.320 70.855 ;
        RECT 51.290 70.585 52.320 70.845 ;
        RECT 51.320 70.405 51.580 70.585 ;
        RECT 51.950 70.575 52.320 70.585 ;
        RECT 53.565 70.405 53.825 71.215 ;
        RECT 58.105 71.205 58.475 71.215 ;
        RECT 57.285 70.845 57.655 70.855 ;
        RECT 56.625 70.585 57.655 70.845 ;
        RECT 56.655 70.405 56.915 70.585 ;
        RECT 57.285 70.575 57.655 70.585 ;
        RECT 58.890 70.405 59.150 71.215 ;
        RECT 63.440 71.205 63.810 71.215 ;
        RECT 62.610 70.845 62.980 70.855 ;
        RECT 61.950 70.585 62.980 70.845 ;
        RECT 61.980 70.405 62.240 70.585 ;
        RECT 62.610 70.575 62.980 70.585 ;
        RECT 64.225 70.405 64.485 71.215 ;
        RECT 68.765 71.205 69.135 71.215 ;
        RECT 67.945 70.845 68.315 70.855 ;
        RECT 67.285 70.585 68.315 70.845 ;
        RECT 67.315 70.405 67.575 70.585 ;
        RECT 67.945 70.575 68.315 70.585 ;
        RECT 69.550 70.405 69.810 71.215 ;
        RECT 74.100 71.205 74.470 71.215 ;
        RECT 73.270 70.845 73.640 70.855 ;
        RECT 72.610 70.585 73.640 70.845 ;
        RECT 72.640 70.405 72.900 70.585 ;
        RECT 73.270 70.575 73.640 70.585 ;
        RECT 74.885 70.405 75.145 71.215 ;
        RECT 79.425 71.205 79.795 71.215 ;
        RECT 78.605 70.845 78.975 70.855 ;
        RECT 77.945 70.585 78.975 70.845 ;
        RECT 77.975 70.405 78.235 70.585 ;
        RECT 78.605 70.575 78.975 70.585 ;
        RECT 80.210 70.405 80.470 71.215 ;
        RECT 84.760 71.205 85.130 71.215 ;
        RECT 83.930 70.845 84.300 70.855 ;
        RECT 83.270 70.585 84.300 70.845 ;
        RECT 83.300 70.405 83.560 70.585 ;
        RECT 83.930 70.575 84.300 70.585 ;
        RECT 85.545 70.405 85.805 71.215 ;
        RECT 90.085 71.205 90.455 71.215 ;
        RECT 89.265 70.845 89.635 70.855 ;
        RECT 88.605 70.585 89.635 70.845 ;
        RECT 88.635 70.405 88.895 70.585 ;
        RECT 89.265 70.575 89.635 70.585 ;
        RECT 90.870 70.405 91.130 71.215 ;
        RECT 95.420 71.205 95.790 71.215 ;
        RECT 94.590 70.845 94.960 70.855 ;
        RECT 93.930 70.585 94.960 70.845 ;
        RECT 93.960 70.405 94.220 70.585 ;
        RECT 94.590 70.575 94.960 70.585 ;
        RECT 96.205 70.405 96.465 71.215 ;
        RECT 100.745 71.205 101.115 71.215 ;
        RECT 99.925 70.845 100.295 70.855 ;
        RECT 99.265 70.585 100.295 70.845 ;
        RECT 99.295 70.405 99.555 70.585 ;
        RECT 99.925 70.575 100.295 70.585 ;
        RECT 101.530 70.405 101.790 71.215 ;
        RECT 106.080 71.205 106.450 71.215 ;
        RECT 105.250 70.845 105.620 70.855 ;
        RECT 104.590 70.585 105.620 70.845 ;
        RECT 104.620 70.405 104.880 70.585 ;
        RECT 105.250 70.575 105.620 70.585 ;
        RECT 106.865 70.405 107.125 71.215 ;
        RECT 111.405 71.205 111.775 71.215 ;
        RECT 110.585 70.845 110.955 70.855 ;
        RECT 109.925 70.585 110.955 70.845 ;
        RECT 109.955 70.405 110.215 70.585 ;
        RECT 110.585 70.575 110.955 70.585 ;
        RECT 112.190 70.405 112.450 71.215 ;
        RECT 116.740 71.205 117.110 71.215 ;
        RECT 115.910 70.845 116.280 70.855 ;
        RECT 115.250 70.585 116.280 70.845 ;
        RECT 115.280 70.405 115.540 70.585 ;
        RECT 115.910 70.575 116.280 70.585 ;
        RECT 117.525 70.405 117.785 71.215 ;
        RECT 122.065 71.205 122.435 71.215 ;
        RECT 121.245 70.845 121.615 70.855 ;
        RECT 120.585 70.585 121.615 70.845 ;
        RECT 120.615 70.405 120.875 70.585 ;
        RECT 121.245 70.575 121.615 70.585 ;
        RECT 122.850 70.405 123.110 71.215 ;
        RECT 126.570 70.845 126.940 70.855 ;
        RECT 125.910 70.585 126.940 70.845 ;
        RECT 125.940 70.405 126.200 70.585 ;
        RECT 126.570 70.575 126.940 70.585 ;
        RECT 127.520 70.405 128.660 76.815 ;
        RECT 31.240 69.280 128.660 70.405 ;
        RECT 31.465 69.110 31.835 69.120 ;
        RECT 32.195 69.110 32.455 69.280 ;
        RECT 31.465 68.850 32.485 69.110 ;
        RECT 31.465 68.840 31.835 68.850 ;
        RECT 35.285 68.460 35.545 69.280 ;
        RECT 74.105 69.110 74.475 69.120 ;
        RECT 116.745 69.110 117.115 69.120 ;
        RECT 122.070 69.110 122.440 69.120 ;
        RECT 122.800 69.110 123.060 69.280 ;
        RECT 74.105 68.850 75.125 69.110 ;
        RECT 116.745 68.850 117.765 69.110 ;
        RECT 122.070 68.850 123.090 69.110 ;
        RECT 74.105 68.840 74.475 68.850 ;
        RECT 116.745 68.840 117.115 68.850 ;
        RECT 122.070 68.840 122.440 68.850 ;
        RECT 35.960 68.460 36.330 68.470 ;
        RECT 125.890 68.460 126.150 69.280 ;
        RECT 126.565 68.460 126.935 68.470 ;
        RECT 35.255 68.200 36.330 68.460 ;
        RECT 125.860 68.200 126.935 68.460 ;
        RECT 35.960 68.190 36.330 68.200 ;
        RECT 126.565 68.190 126.935 68.200 ;
        RECT 31.460 63.940 31.830 63.950 ;
        RECT 122.065 63.940 122.435 63.950 ;
        RECT 31.460 63.680 32.535 63.940 ;
        RECT 122.065 63.680 123.140 63.940 ;
        RECT 31.460 63.670 31.830 63.680 ;
        RECT 32.245 62.870 32.505 63.680 ;
        RECT 122.065 63.670 122.435 63.680 ;
        RECT 35.965 63.310 36.335 63.320 ;
        RECT 35.305 63.050 36.335 63.310 ;
        RECT 35.335 62.870 35.595 63.050 ;
        RECT 35.965 63.040 36.335 63.050 ;
        RECT 122.850 62.870 123.110 63.680 ;
        RECT 126.570 63.310 126.940 63.320 ;
        RECT 125.910 63.050 126.940 63.310 ;
        RECT 125.940 62.870 126.200 63.050 ;
        RECT 126.570 63.040 126.940 63.050 ;
        RECT 127.520 62.870 128.660 69.280 ;
        RECT 31.240 61.745 128.660 62.870 ;
        RECT 31.465 61.575 31.835 61.585 ;
        RECT 32.195 61.575 32.455 61.745 ;
        RECT 31.465 61.315 32.485 61.575 ;
        RECT 31.465 61.305 31.835 61.315 ;
        RECT 35.285 60.925 35.545 61.745 ;
        RECT 122.070 61.575 122.440 61.585 ;
        RECT 122.800 61.575 123.060 61.745 ;
        RECT 122.070 61.315 123.090 61.575 ;
        RECT 122.070 61.305 122.440 61.315 ;
        RECT 35.960 60.925 36.330 60.935 ;
        RECT 125.890 60.925 126.150 61.745 ;
        RECT 126.565 60.925 126.935 60.935 ;
        RECT 35.255 60.665 36.330 60.925 ;
        RECT 125.860 60.665 126.935 60.925 ;
        RECT 35.960 60.655 36.330 60.665 ;
        RECT 126.565 60.655 126.935 60.665 ;
        RECT 31.460 56.405 31.830 56.415 ;
        RECT 122.065 56.405 122.435 56.415 ;
        RECT 31.460 56.145 32.535 56.405 ;
        RECT 122.065 56.145 123.140 56.405 ;
        RECT 31.460 56.135 31.830 56.145 ;
        RECT 32.245 55.335 32.505 56.145 ;
        RECT 122.065 56.135 122.435 56.145 ;
        RECT 35.965 55.775 36.335 55.785 ;
        RECT 35.305 55.515 36.335 55.775 ;
        RECT 35.335 55.335 35.595 55.515 ;
        RECT 35.965 55.505 36.335 55.515 ;
        RECT 122.850 55.335 123.110 56.145 ;
        RECT 126.570 55.775 126.940 55.785 ;
        RECT 125.910 55.515 126.940 55.775 ;
        RECT 125.940 55.335 126.200 55.515 ;
        RECT 126.570 55.505 126.940 55.515 ;
        RECT 127.520 55.335 128.660 61.745 ;
        RECT 31.240 54.210 128.660 55.335 ;
        RECT 31.465 54.040 31.835 54.050 ;
        RECT 32.195 54.040 32.455 54.210 ;
        RECT 31.465 53.780 32.485 54.040 ;
        RECT 31.465 53.770 31.835 53.780 ;
        RECT 35.285 53.390 35.545 54.210 ;
        RECT 122.070 54.040 122.440 54.050 ;
        RECT 122.800 54.040 123.060 54.210 ;
        RECT 122.070 53.780 123.090 54.040 ;
        RECT 122.070 53.770 122.440 53.780 ;
        RECT 35.960 53.390 36.330 53.400 ;
        RECT 125.890 53.390 126.150 54.210 ;
        RECT 126.565 53.390 126.935 53.400 ;
        RECT 35.255 53.130 36.330 53.390 ;
        RECT 125.860 53.130 126.935 53.390 ;
        RECT 35.960 53.120 36.330 53.130 ;
        RECT 126.565 53.120 126.935 53.130 ;
        RECT 31.460 48.870 31.830 48.880 ;
        RECT 122.065 48.870 122.435 48.880 ;
        RECT 31.460 48.610 32.535 48.870 ;
        RECT 122.065 48.610 123.140 48.870 ;
        RECT 31.460 48.600 31.830 48.610 ;
        RECT 32.245 47.800 32.505 48.610 ;
        RECT 122.065 48.600 122.435 48.610 ;
        RECT 35.965 48.240 36.335 48.250 ;
        RECT 35.305 47.980 36.335 48.240 ;
        RECT 35.335 47.800 35.595 47.980 ;
        RECT 35.965 47.970 36.335 47.980 ;
        RECT 122.850 47.800 123.110 48.610 ;
        RECT 126.570 48.240 126.940 48.250 ;
        RECT 125.910 47.980 126.940 48.240 ;
        RECT 125.940 47.800 126.200 47.980 ;
        RECT 126.570 47.970 126.940 47.980 ;
        RECT 127.520 47.800 128.660 54.210 ;
        RECT 31.240 46.675 128.660 47.800 ;
        RECT 31.465 46.505 31.835 46.515 ;
        RECT 32.195 46.505 32.455 46.675 ;
        RECT 31.465 46.245 32.485 46.505 ;
        RECT 31.465 46.235 31.835 46.245 ;
        RECT 35.285 45.855 35.545 46.675 ;
        RECT 122.070 46.505 122.440 46.515 ;
        RECT 122.800 46.505 123.060 46.675 ;
        RECT 122.070 46.245 123.090 46.505 ;
        RECT 122.070 46.235 122.440 46.245 ;
        RECT 35.960 45.855 36.330 45.865 ;
        RECT 125.890 45.855 126.150 46.675 ;
        RECT 126.565 45.855 126.935 45.865 ;
        RECT 35.255 45.595 36.330 45.855 ;
        RECT 125.860 45.595 126.935 45.855 ;
        RECT 35.960 45.585 36.330 45.595 ;
        RECT 126.565 45.585 126.935 45.595 ;
        RECT 31.460 41.335 31.830 41.345 ;
        RECT 122.065 41.335 122.435 41.345 ;
        RECT 31.460 41.075 32.535 41.335 ;
        RECT 122.065 41.075 123.140 41.335 ;
        RECT 31.460 41.065 31.830 41.075 ;
        RECT 32.245 40.265 32.505 41.075 ;
        RECT 122.065 41.065 122.435 41.075 ;
        RECT 35.965 40.705 36.335 40.715 ;
        RECT 35.305 40.445 36.335 40.705 ;
        RECT 35.335 40.265 35.595 40.445 ;
        RECT 35.965 40.435 36.335 40.445 ;
        RECT 122.850 40.265 123.110 41.075 ;
        RECT 126.570 40.705 126.940 40.715 ;
        RECT 125.910 40.445 126.940 40.705 ;
        RECT 125.940 40.265 126.200 40.445 ;
        RECT 126.570 40.435 126.940 40.445 ;
        RECT 127.520 40.265 128.660 46.675 ;
        RECT 31.240 39.140 128.660 40.265 ;
        RECT 31.465 38.970 31.835 38.980 ;
        RECT 32.195 38.970 32.455 39.140 ;
        RECT 31.465 38.710 32.485 38.970 ;
        RECT 31.465 38.700 31.835 38.710 ;
        RECT 35.285 38.320 35.545 39.140 ;
        RECT 122.070 38.970 122.440 38.980 ;
        RECT 122.800 38.970 123.060 39.140 ;
        RECT 122.070 38.710 123.090 38.970 ;
        RECT 122.070 38.700 122.440 38.710 ;
        RECT 35.960 38.320 36.330 38.330 ;
        RECT 125.890 38.320 126.150 39.140 ;
        RECT 126.565 38.320 126.935 38.330 ;
        RECT 35.255 38.060 36.330 38.320 ;
        RECT 125.860 38.060 126.935 38.320 ;
        RECT 35.960 38.050 36.330 38.060 ;
        RECT 126.565 38.050 126.935 38.060 ;
        RECT 31.460 33.800 31.830 33.810 ;
        RECT 122.065 33.800 122.435 33.810 ;
        RECT 31.460 33.540 32.535 33.800 ;
        RECT 122.065 33.540 123.140 33.800 ;
        RECT 31.460 33.530 31.830 33.540 ;
        RECT 32.245 32.730 32.505 33.540 ;
        RECT 122.065 33.530 122.435 33.540 ;
        RECT 35.965 33.170 36.335 33.180 ;
        RECT 35.305 32.910 36.335 33.170 ;
        RECT 35.335 32.730 35.595 32.910 ;
        RECT 35.965 32.900 36.335 32.910 ;
        RECT 122.850 32.730 123.110 33.540 ;
        RECT 126.570 33.170 126.940 33.180 ;
        RECT 125.910 32.910 126.940 33.170 ;
        RECT 125.940 32.730 126.200 32.910 ;
        RECT 126.570 32.900 126.940 32.910 ;
        RECT 127.520 32.730 128.660 39.140 ;
        RECT 31.240 31.605 128.660 32.730 ;
        RECT 31.465 31.435 31.835 31.445 ;
        RECT 32.195 31.435 32.455 31.605 ;
        RECT 31.465 31.175 32.485 31.435 ;
        RECT 31.465 31.165 31.835 31.175 ;
        RECT 35.285 30.785 35.545 31.605 ;
        RECT 122.070 31.435 122.440 31.445 ;
        RECT 122.800 31.435 123.060 31.605 ;
        RECT 122.070 31.175 123.090 31.435 ;
        RECT 122.070 31.165 122.440 31.175 ;
        RECT 35.960 30.785 36.330 30.795 ;
        RECT 125.890 30.785 126.150 31.605 ;
        RECT 126.565 30.785 126.935 30.795 ;
        RECT 35.255 30.525 36.330 30.785 ;
        RECT 125.860 30.525 126.935 30.785 ;
        RECT 35.960 30.515 36.330 30.525 ;
        RECT 126.565 30.515 126.935 30.525 ;
        RECT 31.460 26.265 31.830 26.275 ;
        RECT 122.065 26.265 122.435 26.275 ;
        RECT 31.460 26.005 32.535 26.265 ;
        RECT 122.065 26.005 123.140 26.265 ;
        RECT 31.460 25.995 31.830 26.005 ;
        RECT 32.245 25.195 32.505 26.005 ;
        RECT 122.065 25.995 122.435 26.005 ;
        RECT 35.965 25.635 36.335 25.645 ;
        RECT 35.305 25.375 36.335 25.635 ;
        RECT 35.335 25.195 35.595 25.375 ;
        RECT 35.965 25.365 36.335 25.375 ;
        RECT 122.850 25.195 123.110 26.005 ;
        RECT 126.570 25.635 126.940 25.645 ;
        RECT 125.910 25.375 126.940 25.635 ;
        RECT 125.940 25.195 126.200 25.375 ;
        RECT 126.570 25.365 126.940 25.375 ;
        RECT 127.520 25.195 128.660 31.605 ;
        RECT 31.240 24.070 128.660 25.195 ;
        RECT 31.465 23.900 31.835 23.910 ;
        RECT 32.195 23.900 32.455 24.070 ;
        RECT 31.465 23.640 32.485 23.900 ;
        RECT 31.465 23.630 31.835 23.640 ;
        RECT 35.285 23.250 35.545 24.070 ;
        RECT 122.070 23.900 122.440 23.910 ;
        RECT 122.800 23.900 123.060 24.070 ;
        RECT 122.070 23.640 123.090 23.900 ;
        RECT 122.070 23.630 122.440 23.640 ;
        RECT 35.960 23.250 36.330 23.260 ;
        RECT 125.890 23.250 126.150 24.070 ;
        RECT 126.565 23.250 126.935 23.260 ;
        RECT 35.255 22.990 36.330 23.250 ;
        RECT 125.860 22.990 126.935 23.250 ;
        RECT 35.960 22.980 36.330 22.990 ;
        RECT 126.565 22.980 126.935 22.990 ;
        RECT 31.460 18.730 31.830 18.740 ;
        RECT 122.065 18.730 122.435 18.740 ;
        RECT 31.460 18.470 32.535 18.730 ;
        RECT 122.065 18.470 123.140 18.730 ;
        RECT 31.460 18.460 31.830 18.470 ;
        RECT 32.245 17.660 32.505 18.470 ;
        RECT 122.065 18.460 122.435 18.470 ;
        RECT 35.965 18.100 36.335 18.110 ;
        RECT 35.305 17.840 36.335 18.100 ;
        RECT 35.335 17.660 35.595 17.840 ;
        RECT 35.965 17.830 36.335 17.840 ;
        RECT 122.850 17.660 123.110 18.470 ;
        RECT 126.570 18.100 126.940 18.110 ;
        RECT 125.910 17.840 126.940 18.100 ;
        RECT 125.940 17.660 126.200 17.840 ;
        RECT 126.570 17.830 126.940 17.840 ;
        RECT 127.520 17.660 128.660 24.070 ;
        RECT 31.240 16.535 128.660 17.660 ;
        RECT 31.465 16.365 31.835 16.375 ;
        RECT 32.195 16.365 32.455 16.535 ;
        RECT 31.465 16.105 32.485 16.365 ;
        RECT 31.465 16.095 31.835 16.105 ;
        RECT 35.285 15.715 35.545 16.535 ;
        RECT 122.070 16.365 122.440 16.375 ;
        RECT 122.800 16.365 123.060 16.535 ;
        RECT 122.070 16.105 123.090 16.365 ;
        RECT 122.070 16.095 122.440 16.105 ;
        RECT 35.960 15.715 36.330 15.725 ;
        RECT 125.890 15.715 126.150 16.535 ;
        RECT 126.565 15.715 126.935 15.725 ;
        RECT 35.255 15.455 36.330 15.715 ;
        RECT 125.860 15.455 126.935 15.715 ;
        RECT 35.960 15.445 36.330 15.455 ;
        RECT 126.565 15.445 126.935 15.455 ;
        RECT 31.460 11.195 31.830 11.205 ;
        RECT 122.065 11.195 122.435 11.205 ;
        RECT 31.460 10.935 32.535 11.195 ;
        RECT 122.065 10.935 123.140 11.195 ;
        RECT 31.460 10.925 31.830 10.935 ;
        RECT 32.245 10.125 32.505 10.935 ;
        RECT 122.065 10.925 122.435 10.935 ;
        RECT 35.965 10.565 36.335 10.575 ;
        RECT 35.305 10.305 36.335 10.565 ;
        RECT 35.335 10.125 35.595 10.305 ;
        RECT 35.965 10.295 36.335 10.305 ;
        RECT 122.850 10.125 123.110 10.935 ;
        RECT 126.570 10.565 126.940 10.575 ;
        RECT 125.910 10.305 126.940 10.565 ;
        RECT 125.940 10.125 126.200 10.305 ;
        RECT 126.570 10.295 126.940 10.305 ;
        RECT 127.520 10.125 128.660 16.535 ;
        RECT 31.240 9.000 128.660 10.125 ;
        RECT 31.465 8.830 31.835 8.840 ;
        RECT 32.195 8.830 32.455 9.000 ;
        RECT 31.465 8.570 32.485 8.830 ;
        RECT 31.465 8.560 31.835 8.570 ;
        RECT 35.285 8.180 35.545 9.000 ;
        RECT 36.790 8.830 37.160 8.840 ;
        RECT 37.520 8.830 37.780 9.000 ;
        RECT 36.790 8.570 37.810 8.830 ;
        RECT 36.790 8.560 37.160 8.570 ;
        RECT 35.960 8.180 36.330 8.190 ;
        RECT 40.610 8.180 40.870 9.000 ;
        RECT 42.125 8.830 42.495 8.840 ;
        RECT 42.855 8.830 43.115 9.000 ;
        RECT 42.125 8.570 43.145 8.830 ;
        RECT 42.125 8.560 42.495 8.570 ;
        RECT 41.285 8.180 41.655 8.190 ;
        RECT 45.945 8.180 46.205 9.000 ;
        RECT 47.450 8.830 47.820 8.840 ;
        RECT 48.180 8.830 48.440 9.000 ;
        RECT 47.450 8.570 48.470 8.830 ;
        RECT 47.450 8.560 47.820 8.570 ;
        RECT 46.620 8.180 46.990 8.190 ;
        RECT 51.270 8.180 51.530 9.000 ;
        RECT 52.785 8.830 53.155 8.840 ;
        RECT 53.515 8.830 53.775 9.000 ;
        RECT 52.785 8.570 53.805 8.830 ;
        RECT 52.785 8.560 53.155 8.570 ;
        RECT 51.945 8.180 52.315 8.190 ;
        RECT 56.605 8.180 56.865 9.000 ;
        RECT 58.110 8.830 58.480 8.840 ;
        RECT 58.840 8.830 59.100 9.000 ;
        RECT 58.110 8.570 59.130 8.830 ;
        RECT 58.110 8.560 58.480 8.570 ;
        RECT 57.280 8.180 57.650 8.190 ;
        RECT 61.930 8.180 62.190 9.000 ;
        RECT 63.445 8.830 63.815 8.840 ;
        RECT 64.175 8.830 64.435 9.000 ;
        RECT 63.445 8.570 64.465 8.830 ;
        RECT 63.445 8.560 63.815 8.570 ;
        RECT 62.605 8.180 62.975 8.190 ;
        RECT 67.265 8.180 67.525 9.000 ;
        RECT 68.770 8.830 69.140 8.840 ;
        RECT 69.500 8.830 69.760 9.000 ;
        RECT 68.770 8.570 69.790 8.830 ;
        RECT 68.770 8.560 69.140 8.570 ;
        RECT 67.940 8.180 68.310 8.190 ;
        RECT 72.590 8.180 72.850 9.000 ;
        RECT 74.105 8.830 74.475 8.840 ;
        RECT 74.835 8.830 75.095 9.000 ;
        RECT 74.105 8.570 75.125 8.830 ;
        RECT 74.105 8.560 74.475 8.570 ;
        RECT 73.265 8.180 73.635 8.190 ;
        RECT 77.925 8.180 78.185 9.000 ;
        RECT 79.430 8.830 79.800 8.840 ;
        RECT 80.160 8.830 80.420 9.000 ;
        RECT 79.430 8.570 80.450 8.830 ;
        RECT 79.430 8.560 79.800 8.570 ;
        RECT 78.600 8.180 78.970 8.190 ;
        RECT 83.250 8.180 83.510 9.000 ;
        RECT 84.765 8.830 85.135 8.840 ;
        RECT 85.495 8.830 85.755 9.000 ;
        RECT 84.765 8.570 85.785 8.830 ;
        RECT 84.765 8.560 85.135 8.570 ;
        RECT 83.925 8.180 84.295 8.190 ;
        RECT 88.585 8.180 88.845 9.000 ;
        RECT 90.090 8.830 90.460 8.840 ;
        RECT 90.820 8.830 91.080 9.000 ;
        RECT 90.090 8.570 91.110 8.830 ;
        RECT 90.090 8.560 90.460 8.570 ;
        RECT 89.260 8.180 89.630 8.190 ;
        RECT 93.910 8.180 94.170 9.000 ;
        RECT 95.425 8.830 95.795 8.840 ;
        RECT 96.155 8.830 96.415 9.000 ;
        RECT 95.425 8.570 96.445 8.830 ;
        RECT 95.425 8.560 95.795 8.570 ;
        RECT 94.585 8.180 94.955 8.190 ;
        RECT 99.245 8.180 99.505 9.000 ;
        RECT 100.750 8.830 101.120 8.840 ;
        RECT 101.480 8.830 101.740 9.000 ;
        RECT 100.750 8.570 101.770 8.830 ;
        RECT 100.750 8.560 101.120 8.570 ;
        RECT 99.920 8.180 100.290 8.190 ;
        RECT 104.570 8.180 104.830 9.000 ;
        RECT 106.085 8.830 106.455 8.840 ;
        RECT 106.815 8.830 107.075 9.000 ;
        RECT 106.085 8.570 107.105 8.830 ;
        RECT 106.085 8.560 106.455 8.570 ;
        RECT 105.245 8.180 105.615 8.190 ;
        RECT 109.905 8.180 110.165 9.000 ;
        RECT 111.410 8.830 111.780 8.840 ;
        RECT 112.140 8.830 112.400 9.000 ;
        RECT 111.410 8.570 112.430 8.830 ;
        RECT 111.410 8.560 111.780 8.570 ;
        RECT 110.580 8.180 110.950 8.190 ;
        RECT 115.230 8.180 115.490 9.000 ;
        RECT 116.745 8.830 117.115 8.840 ;
        RECT 117.475 8.830 117.735 9.000 ;
        RECT 116.745 8.570 117.765 8.830 ;
        RECT 116.745 8.560 117.115 8.570 ;
        RECT 115.905 8.180 116.275 8.190 ;
        RECT 120.565 8.180 120.825 9.000 ;
        RECT 122.070 8.830 122.440 8.840 ;
        RECT 122.800 8.830 123.060 9.000 ;
        RECT 122.070 8.570 123.090 8.830 ;
        RECT 122.070 8.560 122.440 8.570 ;
        RECT 121.240 8.180 121.610 8.190 ;
        RECT 125.890 8.180 126.150 9.000 ;
        RECT 126.565 8.180 126.935 8.190 ;
        RECT 35.255 7.920 36.330 8.180 ;
        RECT 40.580 7.920 41.655 8.180 ;
        RECT 45.915 7.920 46.990 8.180 ;
        RECT 51.240 7.920 52.315 8.180 ;
        RECT 56.575 7.920 57.650 8.180 ;
        RECT 61.900 7.920 62.975 8.180 ;
        RECT 67.235 7.920 68.310 8.180 ;
        RECT 72.560 7.920 73.635 8.180 ;
        RECT 77.895 7.920 78.970 8.180 ;
        RECT 83.220 7.920 84.295 8.180 ;
        RECT 88.555 7.920 89.630 8.180 ;
        RECT 93.880 7.920 94.955 8.180 ;
        RECT 99.215 7.920 100.290 8.180 ;
        RECT 104.540 7.920 105.615 8.180 ;
        RECT 109.875 7.920 110.950 8.180 ;
        RECT 115.200 7.920 116.275 8.180 ;
        RECT 120.535 7.920 121.610 8.180 ;
        RECT 125.860 7.920 126.935 8.180 ;
        RECT 35.960 7.910 36.330 7.920 ;
        RECT 41.285 7.910 41.655 7.920 ;
        RECT 46.620 7.910 46.990 7.920 ;
        RECT 51.945 7.910 52.315 7.920 ;
        RECT 57.280 7.910 57.650 7.920 ;
        RECT 62.605 7.910 62.975 7.920 ;
        RECT 67.940 7.910 68.310 7.920 ;
        RECT 73.265 7.910 73.635 7.920 ;
        RECT 78.600 7.910 78.970 7.920 ;
        RECT 83.925 7.910 84.295 7.920 ;
        RECT 89.260 7.910 89.630 7.920 ;
        RECT 94.585 7.910 94.955 7.920 ;
        RECT 99.920 7.910 100.290 7.920 ;
        RECT 105.245 7.910 105.615 7.920 ;
        RECT 110.580 7.910 110.950 7.920 ;
        RECT 115.905 7.910 116.275 7.920 ;
        RECT 121.240 7.910 121.610 7.920 ;
        RECT 126.565 7.910 126.935 7.920 ;
        RECT 31.460 3.660 31.830 3.670 ;
        RECT 36.785 3.660 37.155 3.670 ;
        RECT 42.120 3.660 42.490 3.670 ;
        RECT 47.445 3.660 47.815 3.670 ;
        RECT 52.780 3.660 53.150 3.670 ;
        RECT 58.105 3.660 58.475 3.670 ;
        RECT 63.440 3.660 63.810 3.670 ;
        RECT 68.765 3.660 69.135 3.670 ;
        RECT 74.100 3.660 74.470 3.670 ;
        RECT 79.425 3.660 79.795 3.670 ;
        RECT 84.760 3.660 85.130 3.670 ;
        RECT 90.085 3.660 90.455 3.670 ;
        RECT 95.420 3.660 95.790 3.670 ;
        RECT 100.745 3.660 101.115 3.670 ;
        RECT 106.080 3.660 106.450 3.670 ;
        RECT 111.405 3.660 111.775 3.670 ;
        RECT 116.740 3.660 117.110 3.670 ;
        RECT 122.065 3.660 122.435 3.670 ;
        RECT 31.460 3.400 32.535 3.660 ;
        RECT 36.785 3.400 37.860 3.660 ;
        RECT 42.120 3.400 43.195 3.660 ;
        RECT 47.445 3.400 48.520 3.660 ;
        RECT 52.780 3.400 53.855 3.660 ;
        RECT 58.105 3.400 59.180 3.660 ;
        RECT 63.440 3.400 64.515 3.660 ;
        RECT 68.765 3.400 69.840 3.660 ;
        RECT 74.100 3.400 75.175 3.660 ;
        RECT 79.425 3.400 80.500 3.660 ;
        RECT 84.760 3.400 85.835 3.660 ;
        RECT 90.085 3.400 91.160 3.660 ;
        RECT 95.420 3.400 96.495 3.660 ;
        RECT 100.745 3.400 101.820 3.660 ;
        RECT 106.080 3.400 107.155 3.660 ;
        RECT 111.405 3.400 112.480 3.660 ;
        RECT 116.740 3.400 117.815 3.660 ;
        RECT 122.065 3.400 123.140 3.660 ;
        RECT 31.460 3.390 31.830 3.400 ;
        RECT 32.245 2.590 32.505 3.400 ;
        RECT 36.785 3.390 37.155 3.400 ;
        RECT 35.965 3.030 36.335 3.040 ;
        RECT 35.305 2.770 36.335 3.030 ;
        RECT 35.335 2.590 35.595 2.770 ;
        RECT 35.965 2.760 36.335 2.770 ;
        RECT 37.570 2.590 37.830 3.400 ;
        RECT 42.120 3.390 42.490 3.400 ;
        RECT 41.290 3.030 41.660 3.040 ;
        RECT 40.630 2.770 41.660 3.030 ;
        RECT 40.660 2.590 40.920 2.770 ;
        RECT 41.290 2.760 41.660 2.770 ;
        RECT 42.905 2.590 43.165 3.400 ;
        RECT 47.445 3.390 47.815 3.400 ;
        RECT 46.625 3.030 46.995 3.040 ;
        RECT 45.965 2.770 46.995 3.030 ;
        RECT 45.995 2.590 46.255 2.770 ;
        RECT 46.625 2.760 46.995 2.770 ;
        RECT 48.230 2.590 48.490 3.400 ;
        RECT 52.780 3.390 53.150 3.400 ;
        RECT 51.950 3.030 52.320 3.040 ;
        RECT 51.290 2.770 52.320 3.030 ;
        RECT 51.320 2.590 51.580 2.770 ;
        RECT 51.950 2.760 52.320 2.770 ;
        RECT 53.565 2.590 53.825 3.400 ;
        RECT 58.105 3.390 58.475 3.400 ;
        RECT 57.285 3.030 57.655 3.040 ;
        RECT 56.625 2.770 57.655 3.030 ;
        RECT 56.655 2.590 56.915 2.770 ;
        RECT 57.285 2.760 57.655 2.770 ;
        RECT 58.890 2.590 59.150 3.400 ;
        RECT 63.440 3.390 63.810 3.400 ;
        RECT 62.610 3.030 62.980 3.040 ;
        RECT 61.950 2.770 62.980 3.030 ;
        RECT 61.980 2.590 62.240 2.770 ;
        RECT 62.610 2.760 62.980 2.770 ;
        RECT 64.225 2.590 64.485 3.400 ;
        RECT 68.765 3.390 69.135 3.400 ;
        RECT 67.945 3.030 68.315 3.040 ;
        RECT 67.285 2.770 68.315 3.030 ;
        RECT 67.315 2.590 67.575 2.770 ;
        RECT 67.945 2.760 68.315 2.770 ;
        RECT 69.550 2.590 69.810 3.400 ;
        RECT 74.100 3.390 74.470 3.400 ;
        RECT 73.270 3.030 73.640 3.040 ;
        RECT 72.610 2.770 73.640 3.030 ;
        RECT 72.640 2.590 72.900 2.770 ;
        RECT 73.270 2.760 73.640 2.770 ;
        RECT 74.885 2.590 75.145 3.400 ;
        RECT 79.425 3.390 79.795 3.400 ;
        RECT 78.605 3.030 78.975 3.040 ;
        RECT 77.945 2.770 78.975 3.030 ;
        RECT 77.975 2.590 78.235 2.770 ;
        RECT 78.605 2.760 78.975 2.770 ;
        RECT 80.210 2.590 80.470 3.400 ;
        RECT 84.760 3.390 85.130 3.400 ;
        RECT 83.930 3.030 84.300 3.040 ;
        RECT 83.270 2.770 84.300 3.030 ;
        RECT 83.300 2.590 83.560 2.770 ;
        RECT 83.930 2.760 84.300 2.770 ;
        RECT 85.545 2.590 85.805 3.400 ;
        RECT 90.085 3.390 90.455 3.400 ;
        RECT 89.265 3.030 89.635 3.040 ;
        RECT 88.605 2.770 89.635 3.030 ;
        RECT 88.635 2.590 88.895 2.770 ;
        RECT 89.265 2.760 89.635 2.770 ;
        RECT 90.870 2.590 91.130 3.400 ;
        RECT 95.420 3.390 95.790 3.400 ;
        RECT 94.590 3.030 94.960 3.040 ;
        RECT 93.930 2.770 94.960 3.030 ;
        RECT 93.960 2.590 94.220 2.770 ;
        RECT 94.590 2.760 94.960 2.770 ;
        RECT 96.205 2.590 96.465 3.400 ;
        RECT 100.745 3.390 101.115 3.400 ;
        RECT 99.925 3.030 100.295 3.040 ;
        RECT 99.265 2.770 100.295 3.030 ;
        RECT 99.295 2.590 99.555 2.770 ;
        RECT 99.925 2.760 100.295 2.770 ;
        RECT 101.530 2.590 101.790 3.400 ;
        RECT 106.080 3.390 106.450 3.400 ;
        RECT 105.250 3.030 105.620 3.040 ;
        RECT 104.590 2.770 105.620 3.030 ;
        RECT 104.620 2.590 104.880 2.770 ;
        RECT 105.250 2.760 105.620 2.770 ;
        RECT 106.865 2.590 107.125 3.400 ;
        RECT 111.405 3.390 111.775 3.400 ;
        RECT 110.585 3.030 110.955 3.040 ;
        RECT 109.925 2.770 110.955 3.030 ;
        RECT 109.955 2.590 110.215 2.770 ;
        RECT 110.585 2.760 110.955 2.770 ;
        RECT 112.190 2.590 112.450 3.400 ;
        RECT 116.740 3.390 117.110 3.400 ;
        RECT 115.910 3.030 116.280 3.040 ;
        RECT 115.250 2.770 116.280 3.030 ;
        RECT 115.280 2.590 115.540 2.770 ;
        RECT 115.910 2.760 116.280 2.770 ;
        RECT 117.525 2.590 117.785 3.400 ;
        RECT 122.065 3.390 122.435 3.400 ;
        RECT 121.245 3.030 121.615 3.040 ;
        RECT 120.585 2.770 121.615 3.030 ;
        RECT 120.615 2.590 120.875 2.770 ;
        RECT 121.245 2.760 121.615 2.770 ;
        RECT 122.850 2.590 123.110 3.400 ;
        RECT 126.570 3.030 126.940 3.040 ;
        RECT 125.910 2.770 126.940 3.030 ;
        RECT 125.940 2.590 126.200 2.770 ;
        RECT 126.570 2.760 126.940 2.770 ;
        RECT 127.520 2.590 128.660 9.000 ;
        RECT 31.240 1.085 128.660 2.590 ;
        RECT 127.520 1.045 128.660 1.085 ;
      LAYER met3 ;
        RECT 125.740 84.500 128.670 84.505 ;
        RECT 74.775 81.125 75.105 81.455 ;
        RECT 78.955 81.310 128.670 84.500 ;
        RECT 31.485 75.955 31.815 76.705 ;
        RECT 35.980 75.305 36.310 76.055 ;
        RECT 36.810 75.955 37.140 76.705 ;
        RECT 41.305 75.305 41.635 76.055 ;
        RECT 42.145 75.955 42.475 76.705 ;
        RECT 46.640 75.305 46.970 76.055 ;
        RECT 47.470 75.955 47.800 76.705 ;
        RECT 51.965 75.305 52.295 76.055 ;
        RECT 52.805 75.955 53.135 76.705 ;
        RECT 57.300 75.305 57.630 76.055 ;
        RECT 58.130 75.955 58.460 76.705 ;
        RECT 62.625 75.305 62.955 76.055 ;
        RECT 63.465 75.955 63.795 76.705 ;
        RECT 67.960 75.305 68.290 76.055 ;
        RECT 68.790 75.955 69.120 76.705 ;
        RECT 73.285 75.305 73.615 76.055 ;
        RECT 74.125 75.955 74.455 76.705 ;
        RECT 18.195 71.820 21.620 75.030 ;
        RECT 18.195 71.540 21.615 71.820 ;
        RECT 4.130 68.200 21.615 71.540 ;
        RECT 31.480 71.155 31.810 71.905 ;
        RECT 35.985 70.525 36.315 71.275 ;
        RECT 36.805 71.155 37.135 71.905 ;
        RECT 41.310 70.525 41.640 71.275 ;
        RECT 42.140 71.155 42.470 71.905 ;
        RECT 46.645 70.525 46.975 71.275 ;
        RECT 47.465 71.155 47.795 71.905 ;
        RECT 51.970 70.525 52.300 71.275 ;
        RECT 52.800 71.155 53.130 71.905 ;
        RECT 57.305 70.525 57.635 71.275 ;
        RECT 58.125 71.155 58.455 71.905 ;
        RECT 62.630 70.525 62.960 71.275 ;
        RECT 63.460 71.155 63.790 71.905 ;
        RECT 67.965 70.525 68.295 71.275 ;
        RECT 68.785 71.155 69.115 71.905 ;
        RECT 73.290 70.525 73.620 71.275 ;
        RECT 74.120 71.155 74.450 71.905 ;
        RECT 74.790 69.820 75.090 81.125 ;
        RECT 78.620 75.305 78.950 76.055 ;
        RECT 79.450 75.955 79.780 76.705 ;
        RECT 83.945 75.305 84.275 76.055 ;
        RECT 84.785 75.955 85.115 76.705 ;
        RECT 89.280 75.305 89.610 76.055 ;
        RECT 90.110 75.955 90.440 76.705 ;
        RECT 94.605 75.305 94.935 76.055 ;
        RECT 95.445 75.955 95.775 76.705 ;
        RECT 99.940 75.305 100.270 76.055 ;
        RECT 100.770 75.955 101.100 76.705 ;
        RECT 105.265 75.305 105.595 76.055 ;
        RECT 106.105 75.955 106.435 76.705 ;
        RECT 110.600 75.305 110.930 76.055 ;
        RECT 111.430 75.955 111.760 76.705 ;
        RECT 115.925 75.305 116.255 76.055 ;
        RECT 116.765 75.955 117.095 76.705 ;
        RECT 78.625 70.525 78.955 71.275 ;
        RECT 79.445 71.155 79.775 71.905 ;
        RECT 83.950 70.525 84.280 71.275 ;
        RECT 84.780 71.155 85.110 71.905 ;
        RECT 89.285 70.525 89.615 71.275 ;
        RECT 90.105 71.155 90.435 71.905 ;
        RECT 94.610 70.525 94.940 71.275 ;
        RECT 95.440 71.155 95.770 71.905 ;
        RECT 99.945 70.525 100.275 71.275 ;
        RECT 100.765 71.155 101.095 71.905 ;
        RECT 105.270 70.525 105.600 71.275 ;
        RECT 106.100 71.155 106.430 71.905 ;
        RECT 110.605 70.525 110.935 71.275 ;
        RECT 111.425 71.155 111.755 71.905 ;
        RECT 115.930 70.525 116.260 71.275 ;
        RECT 116.760 71.155 117.090 71.905 ;
        RECT 117.430 69.820 117.730 81.310 ;
        RECT 121.260 75.305 121.590 76.055 ;
        RECT 122.090 75.955 122.420 76.705 ;
        RECT 126.585 75.305 126.915 76.055 ;
        RECT 121.265 70.525 121.595 71.275 ;
        RECT 122.085 71.155 122.415 71.905 ;
        RECT 126.590 70.525 126.920 71.275 ;
        RECT 74.125 69.520 75.090 69.820 ;
        RECT 116.765 69.520 117.730 69.820 ;
        RECT 31.485 68.420 31.815 69.170 ;
        RECT 74.125 68.795 74.455 69.520 ;
        RECT 116.765 68.795 117.095 69.520 ;
        RECT 35.980 67.770 36.310 68.520 ;
        RECT 122.090 68.420 122.420 69.170 ;
        RECT 126.585 67.770 126.915 68.520 ;
        RECT 31.480 63.620 31.810 64.370 ;
        RECT 35.985 62.990 36.315 63.740 ;
        RECT 122.085 63.620 122.415 64.370 ;
        RECT 126.590 62.990 126.920 63.740 ;
        RECT 31.485 60.885 31.815 61.635 ;
        RECT 35.980 60.235 36.310 60.985 ;
        RECT 122.090 60.885 122.420 61.635 ;
        RECT 126.585 60.235 126.915 60.985 ;
        RECT 31.480 56.085 31.810 56.835 ;
        RECT 35.985 55.455 36.315 56.205 ;
        RECT 122.085 56.085 122.415 56.835 ;
        RECT 126.590 55.455 126.920 56.205 ;
        RECT 31.485 53.350 31.815 54.100 ;
        RECT 35.980 52.700 36.310 53.450 ;
        RECT 122.090 53.350 122.420 54.100 ;
        RECT 126.585 52.700 126.915 53.450 ;
        RECT 31.480 48.550 31.810 49.300 ;
        RECT 35.985 47.920 36.315 48.670 ;
        RECT 122.085 48.550 122.415 49.300 ;
        RECT 126.590 47.920 126.920 48.670 ;
        RECT 31.485 45.815 31.815 46.565 ;
        RECT 35.980 45.165 36.310 45.915 ;
        RECT 122.090 45.815 122.420 46.565 ;
        RECT 126.585 45.165 126.915 45.915 ;
        RECT 31.480 41.015 31.810 41.765 ;
        RECT 35.985 40.385 36.315 41.135 ;
        RECT 122.085 41.015 122.415 41.765 ;
        RECT 126.590 40.385 126.920 41.135 ;
        RECT 31.485 38.280 31.815 39.030 ;
        RECT 35.980 37.630 36.310 38.380 ;
        RECT 122.090 38.280 122.420 39.030 ;
        RECT 126.585 37.630 126.915 38.380 ;
        RECT 31.480 33.480 31.810 34.230 ;
        RECT 35.985 32.850 36.315 33.600 ;
        RECT 122.085 33.480 122.415 34.230 ;
        RECT 126.590 32.850 126.920 33.600 ;
        RECT 31.485 30.745 31.815 31.495 ;
        RECT 35.980 30.095 36.310 30.845 ;
        RECT 122.090 30.745 122.420 31.495 ;
        RECT 126.585 30.095 126.915 30.845 ;
        RECT 31.480 25.945 31.810 26.695 ;
        RECT 35.985 25.315 36.315 26.065 ;
        RECT 122.085 25.945 122.415 26.695 ;
        RECT 126.590 25.315 126.920 26.065 ;
        RECT 31.485 23.210 31.815 23.960 ;
        RECT 35.980 22.560 36.310 23.310 ;
        RECT 122.090 23.210 122.420 23.960 ;
        RECT 126.585 22.560 126.915 23.310 ;
        RECT 31.480 18.410 31.810 19.160 ;
        RECT 35.985 17.780 36.315 18.530 ;
        RECT 122.085 18.410 122.415 19.160 ;
        RECT 126.590 17.780 126.920 18.530 ;
        RECT 31.485 15.675 31.815 16.425 ;
        RECT 35.980 15.025 36.310 15.775 ;
        RECT 122.090 15.675 122.420 16.425 ;
        RECT 126.585 15.025 126.915 15.775 ;
        RECT 31.480 10.875 31.810 11.625 ;
        RECT 35.985 10.245 36.315 10.995 ;
        RECT 122.085 10.875 122.415 11.625 ;
        RECT 126.590 10.245 126.920 10.995 ;
        RECT 31.485 8.140 31.815 8.890 ;
        RECT 35.980 7.490 36.310 8.240 ;
        RECT 36.810 8.140 37.140 8.890 ;
        RECT 41.305 7.490 41.635 8.240 ;
        RECT 42.145 8.140 42.475 8.890 ;
        RECT 46.640 7.490 46.970 8.240 ;
        RECT 47.470 8.140 47.800 8.890 ;
        RECT 51.965 7.490 52.295 8.240 ;
        RECT 52.805 8.140 53.135 8.890 ;
        RECT 57.300 7.490 57.630 8.240 ;
        RECT 58.130 8.140 58.460 8.890 ;
        RECT 62.625 7.490 62.955 8.240 ;
        RECT 63.465 8.140 63.795 8.890 ;
        RECT 67.960 7.490 68.290 8.240 ;
        RECT 68.790 8.140 69.120 8.890 ;
        RECT 73.285 7.490 73.615 8.240 ;
        RECT 74.125 8.140 74.455 8.890 ;
        RECT 78.620 7.490 78.950 8.240 ;
        RECT 79.450 8.140 79.780 8.890 ;
        RECT 83.945 7.490 84.275 8.240 ;
        RECT 84.785 8.140 85.115 8.890 ;
        RECT 89.280 7.490 89.610 8.240 ;
        RECT 90.110 8.140 90.440 8.890 ;
        RECT 94.605 7.490 94.935 8.240 ;
        RECT 95.445 8.140 95.775 8.890 ;
        RECT 99.940 7.490 100.270 8.240 ;
        RECT 100.770 8.140 101.100 8.890 ;
        RECT 105.265 7.490 105.595 8.240 ;
        RECT 106.105 8.140 106.435 8.890 ;
        RECT 110.600 7.490 110.930 8.240 ;
        RECT 111.430 8.140 111.760 8.890 ;
        RECT 115.925 7.490 116.255 8.240 ;
        RECT 116.765 8.140 117.095 8.890 ;
        RECT 121.260 7.490 121.590 8.240 ;
        RECT 122.090 8.140 122.420 8.890 ;
        RECT 126.585 7.490 126.915 8.240 ;
        RECT 31.480 3.340 31.810 4.090 ;
        RECT 32.935 3.010 34.070 3.215 ;
        RECT 27.580 0.910 34.070 3.010 ;
        RECT 35.985 2.710 36.315 3.460 ;
        RECT 36.805 3.340 37.135 4.090 ;
        RECT 41.310 2.710 41.640 3.460 ;
        RECT 42.140 3.340 42.470 4.090 ;
        RECT 46.645 2.710 46.975 3.460 ;
        RECT 47.465 3.340 47.795 4.090 ;
        RECT 51.970 2.710 52.300 3.460 ;
        RECT 52.800 3.340 53.130 4.090 ;
        RECT 57.305 2.710 57.635 3.460 ;
        RECT 58.125 3.340 58.455 4.090 ;
        RECT 62.630 2.710 62.960 3.460 ;
        RECT 63.460 3.340 63.790 4.090 ;
        RECT 67.965 2.710 68.295 3.460 ;
        RECT 68.785 3.340 69.115 4.090 ;
        RECT 73.290 2.710 73.620 3.460 ;
        RECT 74.120 3.340 74.450 4.090 ;
        RECT 78.625 2.710 78.955 3.460 ;
        RECT 79.445 3.340 79.775 4.090 ;
        RECT 83.950 2.710 84.280 3.460 ;
        RECT 84.780 3.340 85.110 4.090 ;
        RECT 89.285 2.710 89.615 3.460 ;
        RECT 90.105 3.340 90.435 4.090 ;
        RECT 94.610 2.710 94.940 3.460 ;
        RECT 95.440 3.340 95.770 4.090 ;
        RECT 99.945 2.710 100.275 3.460 ;
        RECT 100.765 3.340 101.095 4.090 ;
        RECT 105.270 2.710 105.600 3.460 ;
        RECT 106.100 3.340 106.430 4.090 ;
        RECT 110.605 2.710 110.935 3.460 ;
        RECT 111.425 3.340 111.755 4.090 ;
        RECT 115.930 2.710 116.260 3.460 ;
        RECT 116.760 3.340 117.090 4.090 ;
        RECT 121.265 2.710 121.595 3.460 ;
        RECT 122.085 3.340 122.415 4.090 ;
        RECT 126.590 2.710 126.920 3.460 ;
        RECT 31.695 -0.020 34.070 0.910 ;
      LAYER met4 ;
        RECT -1.000 81.400 129.360 84.500 ;
        RECT 18.195 75.000 21.620 81.400 ;
        RECT 31.485 76.360 31.815 76.375 ;
        RECT 36.810 76.360 37.140 76.375 ;
        RECT 42.145 76.360 42.475 76.375 ;
        RECT 47.470 76.360 47.800 76.375 ;
        RECT 52.805 76.360 53.135 76.375 ;
        RECT 58.130 76.360 58.460 76.375 ;
        RECT 63.465 76.360 63.795 76.375 ;
        RECT 68.790 76.360 69.120 76.375 ;
        RECT 74.125 76.360 74.455 76.375 ;
        RECT 79.450 76.360 79.780 76.375 ;
        RECT 84.785 76.360 85.115 76.375 ;
        RECT 90.110 76.360 90.440 76.375 ;
        RECT 95.445 76.360 95.775 76.375 ;
        RECT 100.770 76.360 101.100 76.375 ;
        RECT 106.105 76.360 106.435 76.375 ;
        RECT 111.430 76.360 111.760 76.375 ;
        RECT 116.765 76.360 117.095 76.375 ;
        RECT 122.090 76.360 122.420 76.375 ;
        RECT 31.240 76.060 127.180 76.360 ;
        RECT 31.485 76.045 31.815 76.060 ;
        RECT 36.810 76.045 37.140 76.060 ;
        RECT 42.145 76.045 42.475 76.060 ;
        RECT 47.470 76.045 47.800 76.060 ;
        RECT 52.805 76.045 53.135 76.060 ;
        RECT 58.130 76.045 58.460 76.060 ;
        RECT 63.465 76.045 63.795 76.060 ;
        RECT 68.790 76.045 69.120 76.060 ;
        RECT 74.125 76.045 74.455 76.060 ;
        RECT 79.450 76.045 79.780 76.060 ;
        RECT 84.785 76.045 85.115 76.060 ;
        RECT 90.110 76.045 90.440 76.060 ;
        RECT 95.445 76.045 95.775 76.060 ;
        RECT 100.770 76.045 101.100 76.060 ;
        RECT 106.105 76.045 106.435 76.060 ;
        RECT 111.430 76.045 111.760 76.060 ;
        RECT 116.765 76.045 117.095 76.060 ;
        RECT 122.090 76.045 122.420 76.060 ;
        RECT 35.980 75.715 36.310 75.730 ;
        RECT 41.305 75.715 41.635 75.730 ;
        RECT 46.640 75.715 46.970 75.730 ;
        RECT 51.965 75.715 52.295 75.730 ;
        RECT 57.300 75.715 57.630 75.730 ;
        RECT 62.625 75.715 62.955 75.730 ;
        RECT 67.960 75.715 68.290 75.730 ;
        RECT 73.285 75.715 73.615 75.730 ;
        RECT 78.620 75.715 78.950 75.730 ;
        RECT 83.945 75.715 84.275 75.730 ;
        RECT 89.280 75.715 89.610 75.730 ;
        RECT 94.605 75.715 94.935 75.730 ;
        RECT 99.940 75.715 100.270 75.730 ;
        RECT 105.265 75.715 105.595 75.730 ;
        RECT 110.600 75.715 110.930 75.730 ;
        RECT 115.925 75.715 116.255 75.730 ;
        RECT 121.260 75.715 121.590 75.730 ;
        RECT 126.585 75.715 126.915 75.730 ;
        RECT 31.240 75.415 127.180 75.715 ;
        RECT 35.980 75.400 36.310 75.415 ;
        RECT 41.305 75.400 41.635 75.415 ;
        RECT 46.640 75.400 46.970 75.415 ;
        RECT 51.965 75.400 52.295 75.415 ;
        RECT 57.300 75.400 57.630 75.415 ;
        RECT 62.625 75.400 62.955 75.415 ;
        RECT 67.960 75.400 68.290 75.415 ;
        RECT 73.285 75.400 73.615 75.415 ;
        RECT 78.620 75.400 78.950 75.415 ;
        RECT 83.945 75.400 84.275 75.415 ;
        RECT 89.280 75.400 89.610 75.415 ;
        RECT 94.605 75.400 94.935 75.415 ;
        RECT 99.940 75.400 100.270 75.415 ;
        RECT 105.265 75.400 105.595 75.415 ;
        RECT 110.600 75.400 110.930 75.415 ;
        RECT 115.925 75.400 116.255 75.415 ;
        RECT 121.260 75.400 121.590 75.415 ;
        RECT 126.585 75.400 126.915 75.415 ;
        RECT 18.160 71.900 29.345 75.000 ;
        RECT 27.585 0.330 29.345 71.900 ;
        RECT 31.480 71.800 31.810 71.810 ;
        RECT 36.805 71.800 37.135 71.810 ;
        RECT 42.140 71.800 42.470 71.810 ;
        RECT 47.465 71.800 47.795 71.810 ;
        RECT 52.800 71.800 53.130 71.810 ;
        RECT 58.125 71.800 58.455 71.810 ;
        RECT 63.460 71.800 63.790 71.810 ;
        RECT 68.785 71.800 69.115 71.810 ;
        RECT 74.120 71.800 74.450 71.810 ;
        RECT 79.445 71.800 79.775 71.810 ;
        RECT 84.780 71.800 85.110 71.810 ;
        RECT 90.105 71.800 90.435 71.810 ;
        RECT 95.440 71.800 95.770 71.810 ;
        RECT 100.765 71.800 101.095 71.810 ;
        RECT 106.100 71.800 106.430 71.810 ;
        RECT 111.425 71.800 111.755 71.810 ;
        RECT 116.760 71.800 117.090 71.810 ;
        RECT 122.085 71.800 122.415 71.810 ;
        RECT 31.240 71.500 127.180 71.800 ;
        RECT 31.480 71.480 31.810 71.500 ;
        RECT 36.805 71.480 37.135 71.500 ;
        RECT 42.140 71.480 42.470 71.500 ;
        RECT 47.465 71.480 47.795 71.500 ;
        RECT 52.800 71.480 53.130 71.500 ;
        RECT 58.125 71.480 58.455 71.500 ;
        RECT 63.460 71.480 63.790 71.500 ;
        RECT 68.785 71.480 69.115 71.500 ;
        RECT 74.120 71.480 74.450 71.500 ;
        RECT 79.445 71.480 79.775 71.500 ;
        RECT 84.780 71.480 85.110 71.500 ;
        RECT 90.105 71.480 90.435 71.500 ;
        RECT 95.440 71.480 95.770 71.500 ;
        RECT 100.765 71.480 101.095 71.500 ;
        RECT 106.100 71.480 106.430 71.500 ;
        RECT 111.425 71.480 111.755 71.500 ;
        RECT 116.760 71.480 117.090 71.500 ;
        RECT 122.085 71.480 122.415 71.500 ;
        RECT 35.985 71.155 36.315 71.180 ;
        RECT 41.310 71.155 41.640 71.180 ;
        RECT 46.645 71.155 46.975 71.180 ;
        RECT 51.970 71.155 52.300 71.180 ;
        RECT 57.305 71.155 57.635 71.180 ;
        RECT 62.630 71.155 62.960 71.180 ;
        RECT 67.965 71.155 68.295 71.180 ;
        RECT 73.290 71.155 73.620 71.180 ;
        RECT 78.625 71.155 78.955 71.180 ;
        RECT 83.950 71.155 84.280 71.180 ;
        RECT 89.285 71.155 89.615 71.180 ;
        RECT 94.610 71.155 94.940 71.180 ;
        RECT 99.945 71.155 100.275 71.180 ;
        RECT 105.270 71.155 105.600 71.180 ;
        RECT 110.605 71.155 110.935 71.180 ;
        RECT 115.930 71.155 116.260 71.180 ;
        RECT 121.265 71.155 121.595 71.180 ;
        RECT 126.590 71.155 126.920 71.180 ;
        RECT 31.240 70.855 127.180 71.155 ;
        RECT 35.985 70.850 36.315 70.855 ;
        RECT 41.310 70.850 41.640 70.855 ;
        RECT 46.645 70.850 46.975 70.855 ;
        RECT 51.970 70.850 52.300 70.855 ;
        RECT 57.305 70.850 57.635 70.855 ;
        RECT 62.630 70.850 62.960 70.855 ;
        RECT 67.965 70.850 68.295 70.855 ;
        RECT 73.290 70.850 73.620 70.855 ;
        RECT 78.625 70.850 78.955 70.855 ;
        RECT 83.950 70.850 84.280 70.855 ;
        RECT 89.285 70.850 89.615 70.855 ;
        RECT 94.610 70.850 94.940 70.855 ;
        RECT 99.945 70.850 100.275 70.855 ;
        RECT 105.270 70.850 105.600 70.855 ;
        RECT 110.605 70.850 110.935 70.855 ;
        RECT 115.930 70.850 116.260 70.855 ;
        RECT 121.265 70.850 121.595 70.855 ;
        RECT 126.590 70.850 126.920 70.855 ;
        RECT 31.485 8.545 31.815 8.560 ;
        RECT 36.810 8.545 37.140 8.560 ;
        RECT 42.145 8.545 42.475 8.560 ;
        RECT 47.470 8.545 47.800 8.560 ;
        RECT 52.805 8.545 53.135 8.560 ;
        RECT 58.130 8.545 58.460 8.560 ;
        RECT 63.465 8.545 63.795 8.560 ;
        RECT 68.790 8.545 69.120 8.560 ;
        RECT 74.125 8.545 74.455 8.560 ;
        RECT 79.450 8.545 79.780 8.560 ;
        RECT 84.785 8.545 85.115 8.560 ;
        RECT 90.110 8.545 90.440 8.560 ;
        RECT 95.445 8.545 95.775 8.560 ;
        RECT 100.770 8.545 101.100 8.560 ;
        RECT 106.105 8.545 106.435 8.560 ;
        RECT 111.430 8.545 111.760 8.560 ;
        RECT 116.765 8.545 117.095 8.560 ;
        RECT 122.090 8.545 122.420 8.560 ;
        RECT 31.240 8.245 127.180 8.545 ;
        RECT 31.485 8.230 31.815 8.245 ;
        RECT 36.810 8.230 37.140 8.245 ;
        RECT 42.145 8.230 42.475 8.245 ;
        RECT 47.470 8.230 47.800 8.245 ;
        RECT 52.805 8.230 53.135 8.245 ;
        RECT 58.130 8.230 58.460 8.245 ;
        RECT 63.465 8.230 63.795 8.245 ;
        RECT 68.790 8.230 69.120 8.245 ;
        RECT 74.125 8.230 74.455 8.245 ;
        RECT 79.450 8.230 79.780 8.245 ;
        RECT 84.785 8.230 85.115 8.245 ;
        RECT 90.110 8.230 90.440 8.245 ;
        RECT 95.445 8.230 95.775 8.245 ;
        RECT 100.770 8.230 101.100 8.245 ;
        RECT 106.105 8.230 106.435 8.245 ;
        RECT 111.430 8.230 111.760 8.245 ;
        RECT 116.765 8.230 117.095 8.245 ;
        RECT 122.090 8.230 122.420 8.245 ;
        RECT 35.980 7.900 36.310 7.915 ;
        RECT 41.305 7.900 41.635 7.915 ;
        RECT 46.640 7.900 46.970 7.915 ;
        RECT 51.965 7.900 52.295 7.915 ;
        RECT 57.300 7.900 57.630 7.915 ;
        RECT 62.625 7.900 62.955 7.915 ;
        RECT 67.960 7.900 68.290 7.915 ;
        RECT 73.285 7.900 73.615 7.915 ;
        RECT 78.620 7.900 78.950 7.915 ;
        RECT 83.945 7.900 84.275 7.915 ;
        RECT 89.280 7.900 89.610 7.915 ;
        RECT 94.605 7.900 94.935 7.915 ;
        RECT 99.940 7.900 100.270 7.915 ;
        RECT 105.265 7.900 105.595 7.915 ;
        RECT 110.600 7.900 110.930 7.915 ;
        RECT 115.925 7.900 116.255 7.915 ;
        RECT 121.260 7.900 121.590 7.915 ;
        RECT 126.585 7.900 126.915 7.915 ;
        RECT 31.240 7.600 127.180 7.900 ;
        RECT 35.980 7.585 36.310 7.600 ;
        RECT 41.305 7.585 41.635 7.600 ;
        RECT 46.640 7.585 46.970 7.600 ;
        RECT 51.965 7.585 52.295 7.600 ;
        RECT 57.300 7.585 57.630 7.600 ;
        RECT 62.625 7.585 62.955 7.600 ;
        RECT 67.960 7.585 68.290 7.600 ;
        RECT 73.285 7.585 73.615 7.600 ;
        RECT 78.620 7.585 78.950 7.600 ;
        RECT 83.945 7.585 84.275 7.600 ;
        RECT 89.280 7.585 89.610 7.600 ;
        RECT 94.605 7.585 94.935 7.600 ;
        RECT 99.940 7.585 100.270 7.600 ;
        RECT 105.265 7.585 105.595 7.600 ;
        RECT 110.600 7.585 110.930 7.600 ;
        RECT 115.925 7.585 116.255 7.600 ;
        RECT 121.260 7.585 121.590 7.600 ;
        RECT 126.585 7.585 126.915 7.600 ;
        RECT 31.480 3.985 31.810 3.995 ;
        RECT 36.805 3.985 37.135 3.995 ;
        RECT 42.140 3.985 42.470 3.995 ;
        RECT 47.465 3.985 47.795 3.995 ;
        RECT 52.800 3.985 53.130 3.995 ;
        RECT 58.125 3.985 58.455 3.995 ;
        RECT 63.460 3.985 63.790 3.995 ;
        RECT 68.785 3.985 69.115 3.995 ;
        RECT 74.120 3.985 74.450 3.995 ;
        RECT 79.445 3.985 79.775 3.995 ;
        RECT 84.780 3.985 85.110 3.995 ;
        RECT 90.105 3.985 90.435 3.995 ;
        RECT 95.440 3.985 95.770 3.995 ;
        RECT 100.765 3.985 101.095 3.995 ;
        RECT 106.100 3.985 106.430 3.995 ;
        RECT 111.425 3.985 111.755 3.995 ;
        RECT 116.760 3.985 117.090 3.995 ;
        RECT 122.085 3.985 122.415 3.995 ;
        RECT 31.240 3.685 127.180 3.985 ;
        RECT 31.480 3.665 31.810 3.685 ;
        RECT 36.805 3.665 37.135 3.685 ;
        RECT 42.140 3.665 42.470 3.685 ;
        RECT 47.465 3.665 47.795 3.685 ;
        RECT 52.800 3.665 53.130 3.685 ;
        RECT 58.125 3.665 58.455 3.685 ;
        RECT 63.460 3.665 63.790 3.685 ;
        RECT 68.785 3.665 69.115 3.685 ;
        RECT 74.120 3.665 74.450 3.685 ;
        RECT 79.445 3.665 79.775 3.685 ;
        RECT 84.780 3.665 85.110 3.685 ;
        RECT 90.105 3.665 90.435 3.685 ;
        RECT 95.440 3.665 95.770 3.685 ;
        RECT 100.765 3.665 101.095 3.685 ;
        RECT 106.100 3.665 106.430 3.685 ;
        RECT 111.425 3.665 111.755 3.685 ;
        RECT 116.760 3.665 117.090 3.685 ;
        RECT 122.085 3.665 122.415 3.685 ;
        RECT 35.985 3.340 36.315 3.365 ;
        RECT 41.310 3.340 41.640 3.365 ;
        RECT 46.645 3.340 46.975 3.365 ;
        RECT 51.970 3.340 52.300 3.365 ;
        RECT 57.305 3.340 57.635 3.365 ;
        RECT 62.630 3.340 62.960 3.365 ;
        RECT 67.965 3.340 68.295 3.365 ;
        RECT 73.290 3.340 73.620 3.365 ;
        RECT 78.625 3.340 78.955 3.365 ;
        RECT 83.950 3.340 84.280 3.365 ;
        RECT 89.285 3.340 89.615 3.365 ;
        RECT 94.610 3.340 94.940 3.365 ;
        RECT 99.945 3.340 100.275 3.365 ;
        RECT 105.270 3.340 105.600 3.365 ;
        RECT 110.605 3.340 110.935 3.365 ;
        RECT 115.930 3.340 116.260 3.365 ;
        RECT 121.265 3.340 121.595 3.365 ;
        RECT 126.590 3.340 126.920 3.365 ;
        RECT 31.240 3.040 127.180 3.340 ;
        RECT 35.985 3.035 36.315 3.040 ;
        RECT 41.310 3.035 41.640 3.040 ;
        RECT 46.645 3.035 46.975 3.040 ;
        RECT 51.970 3.035 52.300 3.040 ;
        RECT 57.305 3.035 57.635 3.040 ;
        RECT 62.630 3.035 62.960 3.040 ;
        RECT 67.965 3.035 68.295 3.040 ;
        RECT 73.290 3.035 73.620 3.040 ;
        RECT 78.625 3.035 78.955 3.040 ;
        RECT 83.950 3.035 84.280 3.040 ;
        RECT 89.285 3.035 89.615 3.040 ;
        RECT 94.610 3.035 94.940 3.040 ;
        RECT 99.945 3.035 100.275 3.040 ;
        RECT 105.270 3.035 105.600 3.040 ;
        RECT 110.605 3.035 110.935 3.040 ;
        RECT 115.930 3.035 116.260 3.040 ;
        RECT 121.265 3.035 121.595 3.040 ;
        RECT 126.590 3.035 126.920 3.040 ;
    END
  END vdd
  PIN vss
    ANTENNAGATEAREA 68.250000 ;
    ANTENNADIFFAREA 35.910000 ;
    PORT
      LAYER li1 ;
        RECT 32.955 73.750 33.455 73.920 ;
        RECT 32.955 73.210 33.455 73.380 ;
        RECT 33.740 73.335 34.065 73.795 ;
        RECT 34.335 73.750 34.835 73.920 ;
        RECT 38.280 73.750 38.780 73.920 ;
        RECT 34.335 73.210 34.835 73.380 ;
        RECT 38.280 73.210 38.780 73.380 ;
        RECT 39.065 73.335 39.390 73.795 ;
        RECT 39.660 73.750 40.160 73.920 ;
        RECT 43.615 73.750 44.115 73.920 ;
        RECT 39.660 73.210 40.160 73.380 ;
        RECT 43.615 73.210 44.115 73.380 ;
        RECT 44.400 73.335 44.725 73.795 ;
        RECT 44.995 73.750 45.495 73.920 ;
        RECT 48.940 73.750 49.440 73.920 ;
        RECT 44.995 73.210 45.495 73.380 ;
        RECT 48.940 73.210 49.440 73.380 ;
        RECT 49.725 73.335 50.050 73.795 ;
        RECT 50.320 73.750 50.820 73.920 ;
        RECT 54.275 73.750 54.775 73.920 ;
        RECT 50.320 73.210 50.820 73.380 ;
        RECT 54.275 73.210 54.775 73.380 ;
        RECT 55.060 73.335 55.385 73.795 ;
        RECT 55.655 73.750 56.155 73.920 ;
        RECT 59.600 73.750 60.100 73.920 ;
        RECT 55.655 73.210 56.155 73.380 ;
        RECT 59.600 73.210 60.100 73.380 ;
        RECT 60.385 73.335 60.710 73.795 ;
        RECT 60.980 73.750 61.480 73.920 ;
        RECT 64.935 73.750 65.435 73.920 ;
        RECT 60.980 73.210 61.480 73.380 ;
        RECT 64.935 73.210 65.435 73.380 ;
        RECT 65.720 73.335 66.045 73.795 ;
        RECT 66.315 73.750 66.815 73.920 ;
        RECT 70.260 73.750 70.760 73.920 ;
        RECT 66.315 73.210 66.815 73.380 ;
        RECT 70.260 73.210 70.760 73.380 ;
        RECT 71.045 73.335 71.370 73.795 ;
        RECT 71.640 73.750 72.140 73.920 ;
        RECT 75.595 73.750 76.095 73.920 ;
        RECT 71.640 73.210 72.140 73.380 ;
        RECT 75.595 73.210 76.095 73.380 ;
        RECT 76.380 73.335 76.705 73.795 ;
        RECT 76.975 73.750 77.475 73.920 ;
        RECT 80.920 73.750 81.420 73.920 ;
        RECT 76.975 73.210 77.475 73.380 ;
        RECT 80.920 73.210 81.420 73.380 ;
        RECT 81.705 73.335 82.030 73.795 ;
        RECT 82.300 73.750 82.800 73.920 ;
        RECT 86.255 73.750 86.755 73.920 ;
        RECT 82.300 73.210 82.800 73.380 ;
        RECT 86.255 73.210 86.755 73.380 ;
        RECT 87.040 73.335 87.365 73.795 ;
        RECT 87.635 73.750 88.135 73.920 ;
        RECT 91.580 73.750 92.080 73.920 ;
        RECT 87.635 73.210 88.135 73.380 ;
        RECT 91.580 73.210 92.080 73.380 ;
        RECT 92.365 73.335 92.690 73.795 ;
        RECT 92.960 73.750 93.460 73.920 ;
        RECT 96.915 73.750 97.415 73.920 ;
        RECT 92.960 73.210 93.460 73.380 ;
        RECT 96.915 73.210 97.415 73.380 ;
        RECT 97.700 73.335 98.025 73.795 ;
        RECT 98.295 73.750 98.795 73.920 ;
        RECT 102.240 73.750 102.740 73.920 ;
        RECT 98.295 73.210 98.795 73.380 ;
        RECT 102.240 73.210 102.740 73.380 ;
        RECT 103.025 73.335 103.350 73.795 ;
        RECT 103.620 73.750 104.120 73.920 ;
        RECT 107.575 73.750 108.075 73.920 ;
        RECT 103.620 73.210 104.120 73.380 ;
        RECT 107.575 73.210 108.075 73.380 ;
        RECT 108.360 73.335 108.685 73.795 ;
        RECT 108.955 73.750 109.455 73.920 ;
        RECT 112.900 73.750 113.400 73.920 ;
        RECT 108.955 73.210 109.455 73.380 ;
        RECT 112.900 73.210 113.400 73.380 ;
        RECT 113.685 73.335 114.010 73.795 ;
        RECT 114.280 73.750 114.780 73.920 ;
        RECT 118.235 73.750 118.735 73.920 ;
        RECT 114.280 73.210 114.780 73.380 ;
        RECT 118.235 73.210 118.735 73.380 ;
        RECT 119.020 73.335 119.345 73.795 ;
        RECT 119.615 73.750 120.115 73.920 ;
        RECT 123.560 73.750 124.060 73.920 ;
        RECT 119.615 73.210 120.115 73.380 ;
        RECT 123.560 73.210 124.060 73.380 ;
        RECT 124.345 73.335 124.670 73.795 ;
        RECT 124.940 73.750 125.440 73.920 ;
        RECT 124.940 73.210 125.440 73.380 ;
        RECT 32.955 66.215 33.455 66.385 ;
        RECT 32.955 65.675 33.455 65.845 ;
        RECT 33.740 65.800 34.065 66.260 ;
        RECT 34.335 66.215 34.835 66.385 ;
        RECT 34.335 65.675 34.835 65.845 ;
        RECT 39.065 65.800 39.390 66.260 ;
        RECT 44.400 65.800 44.725 66.260 ;
        RECT 49.725 65.800 50.050 66.260 ;
        RECT 55.060 65.800 55.385 66.260 ;
        RECT 60.385 65.800 60.710 66.260 ;
        RECT 65.720 65.800 66.045 66.260 ;
        RECT 71.045 65.800 71.370 66.260 ;
        RECT 75.595 66.215 76.095 66.385 ;
        RECT 76.380 65.800 76.705 66.260 ;
        RECT 81.705 65.800 82.030 66.260 ;
        RECT 87.040 65.800 87.365 66.260 ;
        RECT 92.365 65.800 92.690 66.260 ;
        RECT 97.700 65.800 98.025 66.260 ;
        RECT 103.025 65.800 103.350 66.260 ;
        RECT 108.360 65.800 108.685 66.260 ;
        RECT 113.685 65.800 114.010 66.260 ;
        RECT 118.235 66.215 118.735 66.385 ;
        RECT 119.020 65.800 119.345 66.260 ;
        RECT 123.560 66.215 124.060 66.385 ;
        RECT 123.560 65.675 124.060 65.845 ;
        RECT 124.345 65.800 124.670 66.260 ;
        RECT 124.940 66.215 125.440 66.385 ;
        RECT 124.940 65.675 125.440 65.845 ;
        RECT 32.955 58.680 33.455 58.850 ;
        RECT 32.955 58.140 33.455 58.310 ;
        RECT 33.740 58.265 34.065 58.725 ;
        RECT 34.335 58.680 34.835 58.850 ;
        RECT 34.335 58.140 34.835 58.310 ;
        RECT 39.065 58.265 39.390 58.725 ;
        RECT 44.400 58.265 44.725 58.725 ;
        RECT 49.725 58.265 50.050 58.725 ;
        RECT 55.060 58.265 55.385 58.725 ;
        RECT 60.385 58.265 60.710 58.725 ;
        RECT 65.720 58.265 66.045 58.725 ;
        RECT 71.045 58.265 71.370 58.725 ;
        RECT 76.380 58.265 76.705 58.725 ;
        RECT 81.705 58.265 82.030 58.725 ;
        RECT 87.040 58.265 87.365 58.725 ;
        RECT 92.365 58.265 92.690 58.725 ;
        RECT 97.700 58.265 98.025 58.725 ;
        RECT 103.025 58.265 103.350 58.725 ;
        RECT 108.360 58.265 108.685 58.725 ;
        RECT 113.685 58.265 114.010 58.725 ;
        RECT 119.020 58.265 119.345 58.725 ;
        RECT 123.560 58.680 124.060 58.850 ;
        RECT 123.560 58.140 124.060 58.310 ;
        RECT 124.345 58.265 124.670 58.725 ;
        RECT 124.940 58.680 125.440 58.850 ;
        RECT 124.940 58.140 125.440 58.310 ;
        RECT 32.955 51.145 33.455 51.315 ;
        RECT 32.955 50.605 33.455 50.775 ;
        RECT 33.740 50.730 34.065 51.190 ;
        RECT 34.335 51.145 34.835 51.315 ;
        RECT 34.335 50.605 34.835 50.775 ;
        RECT 39.065 50.730 39.390 51.190 ;
        RECT 44.400 50.730 44.725 51.190 ;
        RECT 49.725 50.730 50.050 51.190 ;
        RECT 55.060 50.730 55.385 51.190 ;
        RECT 60.385 50.730 60.710 51.190 ;
        RECT 65.720 50.730 66.045 51.190 ;
        RECT 71.045 50.730 71.370 51.190 ;
        RECT 76.380 50.730 76.705 51.190 ;
        RECT 81.705 50.730 82.030 51.190 ;
        RECT 87.040 50.730 87.365 51.190 ;
        RECT 92.365 50.730 92.690 51.190 ;
        RECT 97.700 50.730 98.025 51.190 ;
        RECT 103.025 50.730 103.350 51.190 ;
        RECT 108.360 50.730 108.685 51.190 ;
        RECT 113.685 50.730 114.010 51.190 ;
        RECT 119.020 50.730 119.345 51.190 ;
        RECT 123.560 51.145 124.060 51.315 ;
        RECT 123.560 50.605 124.060 50.775 ;
        RECT 124.345 50.730 124.670 51.190 ;
        RECT 124.940 51.145 125.440 51.315 ;
        RECT 124.940 50.605 125.440 50.775 ;
        RECT 32.955 43.610 33.455 43.780 ;
        RECT 32.955 43.070 33.455 43.240 ;
        RECT 33.740 43.195 34.065 43.655 ;
        RECT 34.335 43.610 34.835 43.780 ;
        RECT 34.335 43.070 34.835 43.240 ;
        RECT 39.065 43.195 39.390 43.655 ;
        RECT 44.400 43.195 44.725 43.655 ;
        RECT 49.725 43.195 50.050 43.655 ;
        RECT 55.060 43.195 55.385 43.655 ;
        RECT 60.385 43.195 60.710 43.655 ;
        RECT 65.720 43.195 66.045 43.655 ;
        RECT 71.045 43.195 71.370 43.655 ;
        RECT 76.380 43.195 76.705 43.655 ;
        RECT 81.705 43.195 82.030 43.655 ;
        RECT 87.040 43.195 87.365 43.655 ;
        RECT 92.365 43.195 92.690 43.655 ;
        RECT 97.700 43.195 98.025 43.655 ;
        RECT 103.025 43.195 103.350 43.655 ;
        RECT 108.360 43.195 108.685 43.655 ;
        RECT 113.685 43.195 114.010 43.655 ;
        RECT 119.020 43.195 119.345 43.655 ;
        RECT 123.560 43.610 124.060 43.780 ;
        RECT 123.560 43.070 124.060 43.240 ;
        RECT 124.345 43.195 124.670 43.655 ;
        RECT 124.940 43.610 125.440 43.780 ;
        RECT 124.940 43.070 125.440 43.240 ;
        RECT 32.955 36.075 33.455 36.245 ;
        RECT 32.955 35.535 33.455 35.705 ;
        RECT 33.740 35.660 34.065 36.120 ;
        RECT 34.335 36.075 34.835 36.245 ;
        RECT 34.335 35.535 34.835 35.705 ;
        RECT 39.065 35.660 39.390 36.120 ;
        RECT 44.400 35.660 44.725 36.120 ;
        RECT 49.725 35.660 50.050 36.120 ;
        RECT 55.060 35.660 55.385 36.120 ;
        RECT 60.385 35.660 60.710 36.120 ;
        RECT 65.720 35.660 66.045 36.120 ;
        RECT 71.045 35.660 71.370 36.120 ;
        RECT 76.380 35.660 76.705 36.120 ;
        RECT 81.705 35.660 82.030 36.120 ;
        RECT 87.040 35.660 87.365 36.120 ;
        RECT 92.365 35.660 92.690 36.120 ;
        RECT 97.700 35.660 98.025 36.120 ;
        RECT 103.025 35.660 103.350 36.120 ;
        RECT 108.360 35.660 108.685 36.120 ;
        RECT 113.685 35.660 114.010 36.120 ;
        RECT 119.020 35.660 119.345 36.120 ;
        RECT 123.560 36.075 124.060 36.245 ;
        RECT 123.560 35.535 124.060 35.705 ;
        RECT 124.345 35.660 124.670 36.120 ;
        RECT 124.940 36.075 125.440 36.245 ;
        RECT 124.940 35.535 125.440 35.705 ;
        RECT 32.955 28.540 33.455 28.710 ;
        RECT 32.955 28.000 33.455 28.170 ;
        RECT 33.740 28.125 34.065 28.585 ;
        RECT 34.335 28.540 34.835 28.710 ;
        RECT 34.335 28.000 34.835 28.170 ;
        RECT 39.065 28.125 39.390 28.585 ;
        RECT 44.400 28.125 44.725 28.585 ;
        RECT 49.725 28.125 50.050 28.585 ;
        RECT 55.060 28.125 55.385 28.585 ;
        RECT 60.385 28.125 60.710 28.585 ;
        RECT 65.720 28.125 66.045 28.585 ;
        RECT 71.045 28.125 71.370 28.585 ;
        RECT 76.380 28.125 76.705 28.585 ;
        RECT 81.705 28.125 82.030 28.585 ;
        RECT 87.040 28.125 87.365 28.585 ;
        RECT 92.365 28.125 92.690 28.585 ;
        RECT 97.700 28.125 98.025 28.585 ;
        RECT 103.025 28.125 103.350 28.585 ;
        RECT 108.360 28.125 108.685 28.585 ;
        RECT 113.685 28.125 114.010 28.585 ;
        RECT 119.020 28.125 119.345 28.585 ;
        RECT 123.560 28.540 124.060 28.710 ;
        RECT 123.560 28.000 124.060 28.170 ;
        RECT 124.345 28.125 124.670 28.585 ;
        RECT 124.940 28.540 125.440 28.710 ;
        RECT 124.940 28.000 125.440 28.170 ;
        RECT 32.955 21.005 33.455 21.175 ;
        RECT 32.955 20.465 33.455 20.635 ;
        RECT 33.740 20.590 34.065 21.050 ;
        RECT 34.335 21.005 34.835 21.175 ;
        RECT 34.335 20.465 34.835 20.635 ;
        RECT 39.065 20.590 39.390 21.050 ;
        RECT 44.400 20.590 44.725 21.050 ;
        RECT 49.725 20.590 50.050 21.050 ;
        RECT 55.060 20.590 55.385 21.050 ;
        RECT 60.385 20.590 60.710 21.050 ;
        RECT 65.720 20.590 66.045 21.050 ;
        RECT 71.045 20.590 71.370 21.050 ;
        RECT 76.380 20.590 76.705 21.050 ;
        RECT 81.705 20.590 82.030 21.050 ;
        RECT 87.040 20.590 87.365 21.050 ;
        RECT 92.365 20.590 92.690 21.050 ;
        RECT 97.700 20.590 98.025 21.050 ;
        RECT 103.025 20.590 103.350 21.050 ;
        RECT 108.360 20.590 108.685 21.050 ;
        RECT 113.685 20.590 114.010 21.050 ;
        RECT 119.020 20.590 119.345 21.050 ;
        RECT 123.560 21.005 124.060 21.175 ;
        RECT 123.560 20.465 124.060 20.635 ;
        RECT 124.345 20.590 124.670 21.050 ;
        RECT 124.940 21.005 125.440 21.175 ;
        RECT 124.940 20.465 125.440 20.635 ;
        RECT 32.955 13.470 33.455 13.640 ;
        RECT 32.955 12.930 33.455 13.100 ;
        RECT 33.740 13.055 34.065 13.515 ;
        RECT 34.335 13.470 34.835 13.640 ;
        RECT 34.335 12.930 34.835 13.100 ;
        RECT 39.065 13.055 39.390 13.515 ;
        RECT 44.400 13.055 44.725 13.515 ;
        RECT 49.725 13.055 50.050 13.515 ;
        RECT 55.060 13.055 55.385 13.515 ;
        RECT 60.385 13.055 60.710 13.515 ;
        RECT 65.720 13.055 66.045 13.515 ;
        RECT 71.045 13.055 71.370 13.515 ;
        RECT 76.380 13.055 76.705 13.515 ;
        RECT 81.705 13.055 82.030 13.515 ;
        RECT 87.040 13.055 87.365 13.515 ;
        RECT 92.365 13.055 92.690 13.515 ;
        RECT 97.700 13.055 98.025 13.515 ;
        RECT 103.025 13.055 103.350 13.515 ;
        RECT 108.360 13.055 108.685 13.515 ;
        RECT 113.685 13.055 114.010 13.515 ;
        RECT 119.020 13.055 119.345 13.515 ;
        RECT 123.560 13.470 124.060 13.640 ;
        RECT 123.560 12.930 124.060 13.100 ;
        RECT 124.345 13.055 124.670 13.515 ;
        RECT 124.940 13.470 125.440 13.640 ;
        RECT 124.940 12.930 125.440 13.100 ;
        RECT 32.955 5.935 33.455 6.105 ;
        RECT 32.955 5.395 33.455 5.565 ;
        RECT 33.740 5.520 34.065 5.980 ;
        RECT 34.335 5.935 34.835 6.105 ;
        RECT 38.280 5.935 38.780 6.105 ;
        RECT 34.335 5.395 34.835 5.565 ;
        RECT 38.280 5.395 38.780 5.565 ;
        RECT 39.065 5.520 39.390 5.980 ;
        RECT 39.660 5.935 40.160 6.105 ;
        RECT 43.615 5.935 44.115 6.105 ;
        RECT 39.660 5.395 40.160 5.565 ;
        RECT 43.615 5.395 44.115 5.565 ;
        RECT 44.400 5.520 44.725 5.980 ;
        RECT 44.995 5.935 45.495 6.105 ;
        RECT 48.940 5.935 49.440 6.105 ;
        RECT 44.995 5.395 45.495 5.565 ;
        RECT 48.940 5.395 49.440 5.565 ;
        RECT 49.725 5.520 50.050 5.980 ;
        RECT 50.320 5.935 50.820 6.105 ;
        RECT 54.275 5.935 54.775 6.105 ;
        RECT 50.320 5.395 50.820 5.565 ;
        RECT 54.275 5.395 54.775 5.565 ;
        RECT 55.060 5.520 55.385 5.980 ;
        RECT 55.655 5.935 56.155 6.105 ;
        RECT 59.600 5.935 60.100 6.105 ;
        RECT 55.655 5.395 56.155 5.565 ;
        RECT 59.600 5.395 60.100 5.565 ;
        RECT 60.385 5.520 60.710 5.980 ;
        RECT 60.980 5.935 61.480 6.105 ;
        RECT 64.935 5.935 65.435 6.105 ;
        RECT 60.980 5.395 61.480 5.565 ;
        RECT 64.935 5.395 65.435 5.565 ;
        RECT 65.720 5.520 66.045 5.980 ;
        RECT 66.315 5.935 66.815 6.105 ;
        RECT 70.260 5.935 70.760 6.105 ;
        RECT 66.315 5.395 66.815 5.565 ;
        RECT 70.260 5.395 70.760 5.565 ;
        RECT 71.045 5.520 71.370 5.980 ;
        RECT 71.640 5.935 72.140 6.105 ;
        RECT 75.595 5.935 76.095 6.105 ;
        RECT 71.640 5.395 72.140 5.565 ;
        RECT 75.595 5.395 76.095 5.565 ;
        RECT 76.380 5.520 76.705 5.980 ;
        RECT 76.975 5.935 77.475 6.105 ;
        RECT 80.920 5.935 81.420 6.105 ;
        RECT 76.975 5.395 77.475 5.565 ;
        RECT 80.920 5.395 81.420 5.565 ;
        RECT 81.705 5.520 82.030 5.980 ;
        RECT 82.300 5.935 82.800 6.105 ;
        RECT 86.255 5.935 86.755 6.105 ;
        RECT 82.300 5.395 82.800 5.565 ;
        RECT 86.255 5.395 86.755 5.565 ;
        RECT 87.040 5.520 87.365 5.980 ;
        RECT 87.635 5.935 88.135 6.105 ;
        RECT 91.580 5.935 92.080 6.105 ;
        RECT 87.635 5.395 88.135 5.565 ;
        RECT 91.580 5.395 92.080 5.565 ;
        RECT 92.365 5.520 92.690 5.980 ;
        RECT 92.960 5.935 93.460 6.105 ;
        RECT 96.915 5.935 97.415 6.105 ;
        RECT 92.960 5.395 93.460 5.565 ;
        RECT 96.915 5.395 97.415 5.565 ;
        RECT 97.700 5.520 98.025 5.980 ;
        RECT 98.295 5.935 98.795 6.105 ;
        RECT 102.240 5.935 102.740 6.105 ;
        RECT 98.295 5.395 98.795 5.565 ;
        RECT 102.240 5.395 102.740 5.565 ;
        RECT 103.025 5.520 103.350 5.980 ;
        RECT 103.620 5.935 104.120 6.105 ;
        RECT 107.575 5.935 108.075 6.105 ;
        RECT 103.620 5.395 104.120 5.565 ;
        RECT 107.575 5.395 108.075 5.565 ;
        RECT 108.360 5.520 108.685 5.980 ;
        RECT 108.955 5.935 109.455 6.105 ;
        RECT 112.900 5.935 113.400 6.105 ;
        RECT 108.955 5.395 109.455 5.565 ;
        RECT 112.900 5.395 113.400 5.565 ;
        RECT 113.685 5.520 114.010 5.980 ;
        RECT 114.280 5.935 114.780 6.105 ;
        RECT 118.235 5.935 118.735 6.105 ;
        RECT 114.280 5.395 114.780 5.565 ;
        RECT 118.235 5.395 118.735 5.565 ;
        RECT 119.020 5.520 119.345 5.980 ;
        RECT 119.615 5.935 120.115 6.105 ;
        RECT 123.560 5.935 124.060 6.105 ;
        RECT 119.615 5.395 120.115 5.565 ;
        RECT 123.560 5.395 124.060 5.565 ;
        RECT 124.345 5.520 124.670 5.980 ;
        RECT 124.940 5.935 125.440 6.105 ;
        RECT 124.940 5.395 125.440 5.565 ;
      LAYER met1 ;
        RECT 29.785 1.085 30.925 78.295 ;
        RECT 32.195 73.950 32.455 74.830 ;
        RECT 35.335 73.950 35.595 74.740 ;
        RECT 32.195 73.720 33.435 73.950 ;
        RECT 33.765 73.775 34.040 73.840 ;
        RECT 32.195 73.180 33.435 73.410 ;
        RECT 33.710 73.355 34.100 73.775 ;
        RECT 34.355 73.720 35.595 73.950 ;
        RECT 37.520 73.950 37.780 74.830 ;
        RECT 40.660 73.950 40.920 74.740 ;
        RECT 37.520 73.720 38.760 73.950 ;
        RECT 39.090 73.775 39.365 73.840 ;
        RECT 33.765 73.295 34.040 73.355 ;
        RECT 34.355 73.180 35.595 73.410 ;
        RECT 32.195 72.485 32.455 73.180 ;
        RECT 35.335 72.390 35.595 73.180 ;
        RECT 37.520 73.180 38.760 73.410 ;
        RECT 39.035 73.355 39.425 73.775 ;
        RECT 39.680 73.720 40.920 73.950 ;
        RECT 42.855 73.950 43.115 74.830 ;
        RECT 45.995 73.950 46.255 74.740 ;
        RECT 42.855 73.720 44.095 73.950 ;
        RECT 44.425 73.775 44.700 73.840 ;
        RECT 39.090 73.295 39.365 73.355 ;
        RECT 39.680 73.180 40.920 73.410 ;
        RECT 37.520 72.485 37.780 73.180 ;
        RECT 40.660 72.390 40.920 73.180 ;
        RECT 42.855 73.180 44.095 73.410 ;
        RECT 44.370 73.355 44.760 73.775 ;
        RECT 45.015 73.720 46.255 73.950 ;
        RECT 48.180 73.950 48.440 74.830 ;
        RECT 51.320 73.950 51.580 74.740 ;
        RECT 48.180 73.720 49.420 73.950 ;
        RECT 49.750 73.775 50.025 73.840 ;
        RECT 44.425 73.295 44.700 73.355 ;
        RECT 45.015 73.180 46.255 73.410 ;
        RECT 42.855 72.485 43.115 73.180 ;
        RECT 45.995 72.390 46.255 73.180 ;
        RECT 48.180 73.180 49.420 73.410 ;
        RECT 49.695 73.355 50.085 73.775 ;
        RECT 50.340 73.720 51.580 73.950 ;
        RECT 53.515 73.950 53.775 74.830 ;
        RECT 56.655 73.950 56.915 74.740 ;
        RECT 53.515 73.720 54.755 73.950 ;
        RECT 55.085 73.775 55.360 73.840 ;
        RECT 49.750 73.295 50.025 73.355 ;
        RECT 50.340 73.180 51.580 73.410 ;
        RECT 48.180 72.485 48.440 73.180 ;
        RECT 51.320 72.390 51.580 73.180 ;
        RECT 53.515 73.180 54.755 73.410 ;
        RECT 55.030 73.355 55.420 73.775 ;
        RECT 55.675 73.720 56.915 73.950 ;
        RECT 58.840 73.950 59.100 74.830 ;
        RECT 61.980 73.950 62.240 74.740 ;
        RECT 58.840 73.720 60.080 73.950 ;
        RECT 60.410 73.775 60.685 73.840 ;
        RECT 55.085 73.295 55.360 73.355 ;
        RECT 55.675 73.180 56.915 73.410 ;
        RECT 53.515 72.485 53.775 73.180 ;
        RECT 56.655 72.390 56.915 73.180 ;
        RECT 58.840 73.180 60.080 73.410 ;
        RECT 60.355 73.355 60.745 73.775 ;
        RECT 61.000 73.720 62.240 73.950 ;
        RECT 64.175 73.950 64.435 74.830 ;
        RECT 67.315 73.950 67.575 74.740 ;
        RECT 64.175 73.720 65.415 73.950 ;
        RECT 65.745 73.775 66.020 73.840 ;
        RECT 60.410 73.295 60.685 73.355 ;
        RECT 61.000 73.180 62.240 73.410 ;
        RECT 58.840 72.485 59.100 73.180 ;
        RECT 61.980 72.390 62.240 73.180 ;
        RECT 64.175 73.180 65.415 73.410 ;
        RECT 65.690 73.355 66.080 73.775 ;
        RECT 66.335 73.720 67.575 73.950 ;
        RECT 69.500 73.950 69.760 74.830 ;
        RECT 72.640 73.950 72.900 74.740 ;
        RECT 69.500 73.720 70.740 73.950 ;
        RECT 71.070 73.775 71.345 73.840 ;
        RECT 65.745 73.295 66.020 73.355 ;
        RECT 66.335 73.180 67.575 73.410 ;
        RECT 64.175 72.485 64.435 73.180 ;
        RECT 67.315 72.390 67.575 73.180 ;
        RECT 69.500 73.180 70.740 73.410 ;
        RECT 71.015 73.355 71.405 73.775 ;
        RECT 71.660 73.720 72.900 73.950 ;
        RECT 74.835 73.950 75.095 74.830 ;
        RECT 77.975 73.950 78.235 74.740 ;
        RECT 74.835 73.720 76.075 73.950 ;
        RECT 76.405 73.775 76.680 73.840 ;
        RECT 71.070 73.295 71.345 73.355 ;
        RECT 71.660 73.180 72.900 73.410 ;
        RECT 69.500 72.485 69.760 73.180 ;
        RECT 72.640 72.390 72.900 73.180 ;
        RECT 74.835 73.180 76.075 73.410 ;
        RECT 76.350 73.355 76.740 73.775 ;
        RECT 76.995 73.720 78.235 73.950 ;
        RECT 80.160 73.950 80.420 74.830 ;
        RECT 83.300 73.950 83.560 74.740 ;
        RECT 80.160 73.720 81.400 73.950 ;
        RECT 81.730 73.775 82.005 73.840 ;
        RECT 76.405 73.295 76.680 73.355 ;
        RECT 76.995 73.180 78.235 73.410 ;
        RECT 74.835 72.485 75.095 73.180 ;
        RECT 77.975 72.390 78.235 73.180 ;
        RECT 80.160 73.180 81.400 73.410 ;
        RECT 81.675 73.355 82.065 73.775 ;
        RECT 82.320 73.720 83.560 73.950 ;
        RECT 85.495 73.950 85.755 74.830 ;
        RECT 88.635 73.950 88.895 74.740 ;
        RECT 85.495 73.720 86.735 73.950 ;
        RECT 87.065 73.775 87.340 73.840 ;
        RECT 81.730 73.295 82.005 73.355 ;
        RECT 82.320 73.180 83.560 73.410 ;
        RECT 80.160 72.485 80.420 73.180 ;
        RECT 83.300 72.390 83.560 73.180 ;
        RECT 85.495 73.180 86.735 73.410 ;
        RECT 87.010 73.355 87.400 73.775 ;
        RECT 87.655 73.720 88.895 73.950 ;
        RECT 90.820 73.950 91.080 74.830 ;
        RECT 93.960 73.950 94.220 74.740 ;
        RECT 90.820 73.720 92.060 73.950 ;
        RECT 92.390 73.775 92.665 73.840 ;
        RECT 87.065 73.295 87.340 73.355 ;
        RECT 87.655 73.180 88.895 73.410 ;
        RECT 85.495 72.485 85.755 73.180 ;
        RECT 88.635 72.390 88.895 73.180 ;
        RECT 90.820 73.180 92.060 73.410 ;
        RECT 92.335 73.355 92.725 73.775 ;
        RECT 92.980 73.720 94.220 73.950 ;
        RECT 96.155 73.950 96.415 74.830 ;
        RECT 99.295 73.950 99.555 74.740 ;
        RECT 96.155 73.720 97.395 73.950 ;
        RECT 97.725 73.775 98.000 73.840 ;
        RECT 92.390 73.295 92.665 73.355 ;
        RECT 92.980 73.180 94.220 73.410 ;
        RECT 90.820 72.485 91.080 73.180 ;
        RECT 93.960 72.390 94.220 73.180 ;
        RECT 96.155 73.180 97.395 73.410 ;
        RECT 97.670 73.355 98.060 73.775 ;
        RECT 98.315 73.720 99.555 73.950 ;
        RECT 101.480 73.950 101.740 74.830 ;
        RECT 104.620 73.950 104.880 74.740 ;
        RECT 101.480 73.720 102.720 73.950 ;
        RECT 103.050 73.775 103.325 73.840 ;
        RECT 97.725 73.295 98.000 73.355 ;
        RECT 98.315 73.180 99.555 73.410 ;
        RECT 96.155 72.485 96.415 73.180 ;
        RECT 99.295 72.390 99.555 73.180 ;
        RECT 101.480 73.180 102.720 73.410 ;
        RECT 102.995 73.355 103.385 73.775 ;
        RECT 103.640 73.720 104.880 73.950 ;
        RECT 106.815 73.950 107.075 74.830 ;
        RECT 109.955 73.950 110.215 74.740 ;
        RECT 106.815 73.720 108.055 73.950 ;
        RECT 108.385 73.775 108.660 73.840 ;
        RECT 103.050 73.295 103.325 73.355 ;
        RECT 103.640 73.180 104.880 73.410 ;
        RECT 101.480 72.485 101.740 73.180 ;
        RECT 104.620 72.390 104.880 73.180 ;
        RECT 106.815 73.180 108.055 73.410 ;
        RECT 108.330 73.355 108.720 73.775 ;
        RECT 108.975 73.720 110.215 73.950 ;
        RECT 112.140 73.950 112.400 74.830 ;
        RECT 115.280 73.950 115.540 74.740 ;
        RECT 112.140 73.720 113.380 73.950 ;
        RECT 113.710 73.775 113.985 73.840 ;
        RECT 108.385 73.295 108.660 73.355 ;
        RECT 108.975 73.180 110.215 73.410 ;
        RECT 106.815 72.485 107.075 73.180 ;
        RECT 109.955 72.390 110.215 73.180 ;
        RECT 112.140 73.180 113.380 73.410 ;
        RECT 113.655 73.355 114.045 73.775 ;
        RECT 114.300 73.720 115.540 73.950 ;
        RECT 117.475 73.950 117.735 74.830 ;
        RECT 120.615 73.950 120.875 74.740 ;
        RECT 117.475 73.720 118.715 73.950 ;
        RECT 119.045 73.775 119.320 73.840 ;
        RECT 113.710 73.295 113.985 73.355 ;
        RECT 114.300 73.180 115.540 73.410 ;
        RECT 112.140 72.485 112.400 73.180 ;
        RECT 115.280 72.390 115.540 73.180 ;
        RECT 117.475 73.180 118.715 73.410 ;
        RECT 118.990 73.355 119.380 73.775 ;
        RECT 119.635 73.720 120.875 73.950 ;
        RECT 122.800 73.950 123.060 74.830 ;
        RECT 125.940 73.950 126.200 74.740 ;
        RECT 122.800 73.720 124.040 73.950 ;
        RECT 124.370 73.775 124.645 73.840 ;
        RECT 119.045 73.295 119.320 73.355 ;
        RECT 119.635 73.180 120.875 73.410 ;
        RECT 117.475 72.485 117.735 73.180 ;
        RECT 120.615 72.390 120.875 73.180 ;
        RECT 122.800 73.180 124.040 73.410 ;
        RECT 124.315 73.355 124.705 73.775 ;
        RECT 124.960 73.720 126.200 73.950 ;
        RECT 124.370 73.295 124.645 73.355 ;
        RECT 124.960 73.180 126.200 73.410 ;
        RECT 122.800 72.485 123.060 73.180 ;
        RECT 125.940 72.390 126.200 73.180 ;
        RECT 32.195 66.415 32.455 67.295 ;
        RECT 35.335 66.415 35.595 67.205 ;
        RECT 32.195 66.185 33.435 66.415 ;
        RECT 33.765 66.240 34.040 66.305 ;
        RECT 32.195 65.645 33.435 65.875 ;
        RECT 33.710 65.820 34.100 66.240 ;
        RECT 34.355 66.185 35.595 66.415 ;
        RECT 74.835 66.415 75.095 67.295 ;
        RECT 117.475 66.415 117.735 67.295 ;
        RECT 122.800 66.415 123.060 67.295 ;
        RECT 125.940 66.415 126.200 67.205 ;
        RECT 39.090 66.240 39.365 66.305 ;
        RECT 44.425 66.240 44.700 66.305 ;
        RECT 49.750 66.240 50.025 66.305 ;
        RECT 55.085 66.240 55.360 66.305 ;
        RECT 60.410 66.240 60.685 66.305 ;
        RECT 65.745 66.240 66.020 66.305 ;
        RECT 71.070 66.240 71.345 66.305 ;
        RECT 33.765 65.760 34.040 65.820 ;
        RECT 34.355 65.645 35.595 65.875 ;
        RECT 39.035 65.820 39.425 66.240 ;
        RECT 44.370 65.820 44.760 66.240 ;
        RECT 49.695 65.820 50.085 66.240 ;
        RECT 55.030 65.820 55.420 66.240 ;
        RECT 60.355 65.820 60.745 66.240 ;
        RECT 65.690 65.820 66.080 66.240 ;
        RECT 71.015 65.820 71.405 66.240 ;
        RECT 74.835 66.185 76.075 66.415 ;
        RECT 76.405 66.240 76.680 66.305 ;
        RECT 81.730 66.240 82.005 66.305 ;
        RECT 87.065 66.240 87.340 66.305 ;
        RECT 92.390 66.240 92.665 66.305 ;
        RECT 97.725 66.240 98.000 66.305 ;
        RECT 103.050 66.240 103.325 66.305 ;
        RECT 108.385 66.240 108.660 66.305 ;
        RECT 113.710 66.240 113.985 66.305 ;
        RECT 76.350 65.820 76.740 66.240 ;
        RECT 81.675 65.820 82.065 66.240 ;
        RECT 87.010 65.820 87.400 66.240 ;
        RECT 92.335 65.820 92.725 66.240 ;
        RECT 97.670 65.820 98.060 66.240 ;
        RECT 102.995 65.820 103.385 66.240 ;
        RECT 108.330 65.820 108.720 66.240 ;
        RECT 113.655 65.820 114.045 66.240 ;
        RECT 117.475 66.185 118.715 66.415 ;
        RECT 119.045 66.240 119.320 66.305 ;
        RECT 118.990 65.820 119.380 66.240 ;
        RECT 122.800 66.185 124.040 66.415 ;
        RECT 124.370 66.240 124.645 66.305 ;
        RECT 39.090 65.760 39.365 65.820 ;
        RECT 44.425 65.760 44.700 65.820 ;
        RECT 49.750 65.760 50.025 65.820 ;
        RECT 55.085 65.760 55.360 65.820 ;
        RECT 60.410 65.760 60.685 65.820 ;
        RECT 65.745 65.760 66.020 65.820 ;
        RECT 71.070 65.760 71.345 65.820 ;
        RECT 76.405 65.760 76.680 65.820 ;
        RECT 81.730 65.760 82.005 65.820 ;
        RECT 87.065 65.760 87.340 65.820 ;
        RECT 92.390 65.760 92.665 65.820 ;
        RECT 97.725 65.760 98.000 65.820 ;
        RECT 103.050 65.760 103.325 65.820 ;
        RECT 108.385 65.760 108.660 65.820 ;
        RECT 113.710 65.760 113.985 65.820 ;
        RECT 119.045 65.760 119.320 65.820 ;
        RECT 32.195 64.950 32.455 65.645 ;
        RECT 35.335 64.855 35.595 65.645 ;
        RECT 122.800 65.645 124.040 65.875 ;
        RECT 124.315 65.820 124.705 66.240 ;
        RECT 124.960 66.185 126.200 66.415 ;
        RECT 124.370 65.760 124.645 65.820 ;
        RECT 124.960 65.645 126.200 65.875 ;
        RECT 122.800 64.950 123.060 65.645 ;
        RECT 125.940 64.855 126.200 65.645 ;
        RECT 32.195 58.880 32.455 59.760 ;
        RECT 35.335 58.880 35.595 59.670 ;
        RECT 32.195 58.650 33.435 58.880 ;
        RECT 33.765 58.705 34.040 58.770 ;
        RECT 32.195 58.110 33.435 58.340 ;
        RECT 33.710 58.285 34.100 58.705 ;
        RECT 34.355 58.650 35.595 58.880 ;
        RECT 122.800 58.880 123.060 59.760 ;
        RECT 125.940 58.880 126.200 59.670 ;
        RECT 39.090 58.705 39.365 58.770 ;
        RECT 44.425 58.705 44.700 58.770 ;
        RECT 49.750 58.705 50.025 58.770 ;
        RECT 55.085 58.705 55.360 58.770 ;
        RECT 60.410 58.705 60.685 58.770 ;
        RECT 65.745 58.705 66.020 58.770 ;
        RECT 71.070 58.705 71.345 58.770 ;
        RECT 76.405 58.705 76.680 58.770 ;
        RECT 81.730 58.705 82.005 58.770 ;
        RECT 87.065 58.705 87.340 58.770 ;
        RECT 92.390 58.705 92.665 58.770 ;
        RECT 97.725 58.705 98.000 58.770 ;
        RECT 103.050 58.705 103.325 58.770 ;
        RECT 108.385 58.705 108.660 58.770 ;
        RECT 113.710 58.705 113.985 58.770 ;
        RECT 119.045 58.705 119.320 58.770 ;
        RECT 33.765 58.225 34.040 58.285 ;
        RECT 34.355 58.110 35.595 58.340 ;
        RECT 39.035 58.285 39.425 58.705 ;
        RECT 44.370 58.285 44.760 58.705 ;
        RECT 49.695 58.285 50.085 58.705 ;
        RECT 55.030 58.285 55.420 58.705 ;
        RECT 60.355 58.285 60.745 58.705 ;
        RECT 65.690 58.285 66.080 58.705 ;
        RECT 71.015 58.285 71.405 58.705 ;
        RECT 76.350 58.285 76.740 58.705 ;
        RECT 81.675 58.285 82.065 58.705 ;
        RECT 87.010 58.285 87.400 58.705 ;
        RECT 92.335 58.285 92.725 58.705 ;
        RECT 97.670 58.285 98.060 58.705 ;
        RECT 102.995 58.285 103.385 58.705 ;
        RECT 108.330 58.285 108.720 58.705 ;
        RECT 113.655 58.285 114.045 58.705 ;
        RECT 118.990 58.285 119.380 58.705 ;
        RECT 122.800 58.650 124.040 58.880 ;
        RECT 124.370 58.705 124.645 58.770 ;
        RECT 39.090 58.225 39.365 58.285 ;
        RECT 44.425 58.225 44.700 58.285 ;
        RECT 49.750 58.225 50.025 58.285 ;
        RECT 55.085 58.225 55.360 58.285 ;
        RECT 60.410 58.225 60.685 58.285 ;
        RECT 65.745 58.225 66.020 58.285 ;
        RECT 71.070 58.225 71.345 58.285 ;
        RECT 76.405 58.225 76.680 58.285 ;
        RECT 81.730 58.225 82.005 58.285 ;
        RECT 87.065 58.225 87.340 58.285 ;
        RECT 92.390 58.225 92.665 58.285 ;
        RECT 97.725 58.225 98.000 58.285 ;
        RECT 103.050 58.225 103.325 58.285 ;
        RECT 108.385 58.225 108.660 58.285 ;
        RECT 113.710 58.225 113.985 58.285 ;
        RECT 119.045 58.225 119.320 58.285 ;
        RECT 32.195 57.415 32.455 58.110 ;
        RECT 35.335 57.320 35.595 58.110 ;
        RECT 122.800 58.110 124.040 58.340 ;
        RECT 124.315 58.285 124.705 58.705 ;
        RECT 124.960 58.650 126.200 58.880 ;
        RECT 124.370 58.225 124.645 58.285 ;
        RECT 124.960 58.110 126.200 58.340 ;
        RECT 122.800 57.415 123.060 58.110 ;
        RECT 125.940 57.320 126.200 58.110 ;
        RECT 32.195 51.345 32.455 52.225 ;
        RECT 35.335 51.345 35.595 52.135 ;
        RECT 32.195 51.115 33.435 51.345 ;
        RECT 33.765 51.170 34.040 51.235 ;
        RECT 32.195 50.575 33.435 50.805 ;
        RECT 33.710 50.750 34.100 51.170 ;
        RECT 34.355 51.115 35.595 51.345 ;
        RECT 122.800 51.345 123.060 52.225 ;
        RECT 125.940 51.345 126.200 52.135 ;
        RECT 39.090 51.170 39.365 51.235 ;
        RECT 44.425 51.170 44.700 51.235 ;
        RECT 49.750 51.170 50.025 51.235 ;
        RECT 55.085 51.170 55.360 51.235 ;
        RECT 60.410 51.170 60.685 51.235 ;
        RECT 65.745 51.170 66.020 51.235 ;
        RECT 71.070 51.170 71.345 51.235 ;
        RECT 76.405 51.170 76.680 51.235 ;
        RECT 81.730 51.170 82.005 51.235 ;
        RECT 87.065 51.170 87.340 51.235 ;
        RECT 92.390 51.170 92.665 51.235 ;
        RECT 97.725 51.170 98.000 51.235 ;
        RECT 103.050 51.170 103.325 51.235 ;
        RECT 108.385 51.170 108.660 51.235 ;
        RECT 113.710 51.170 113.985 51.235 ;
        RECT 119.045 51.170 119.320 51.235 ;
        RECT 33.765 50.690 34.040 50.750 ;
        RECT 34.355 50.575 35.595 50.805 ;
        RECT 39.035 50.750 39.425 51.170 ;
        RECT 44.370 50.750 44.760 51.170 ;
        RECT 49.695 50.750 50.085 51.170 ;
        RECT 55.030 50.750 55.420 51.170 ;
        RECT 60.355 50.750 60.745 51.170 ;
        RECT 65.690 50.750 66.080 51.170 ;
        RECT 71.015 50.750 71.405 51.170 ;
        RECT 76.350 50.750 76.740 51.170 ;
        RECT 81.675 50.750 82.065 51.170 ;
        RECT 87.010 50.750 87.400 51.170 ;
        RECT 92.335 50.750 92.725 51.170 ;
        RECT 97.670 50.750 98.060 51.170 ;
        RECT 102.995 50.750 103.385 51.170 ;
        RECT 108.330 50.750 108.720 51.170 ;
        RECT 113.655 50.750 114.045 51.170 ;
        RECT 118.990 50.750 119.380 51.170 ;
        RECT 122.800 51.115 124.040 51.345 ;
        RECT 124.370 51.170 124.645 51.235 ;
        RECT 39.090 50.690 39.365 50.750 ;
        RECT 44.425 50.690 44.700 50.750 ;
        RECT 49.750 50.690 50.025 50.750 ;
        RECT 55.085 50.690 55.360 50.750 ;
        RECT 60.410 50.690 60.685 50.750 ;
        RECT 65.745 50.690 66.020 50.750 ;
        RECT 71.070 50.690 71.345 50.750 ;
        RECT 76.405 50.690 76.680 50.750 ;
        RECT 81.730 50.690 82.005 50.750 ;
        RECT 87.065 50.690 87.340 50.750 ;
        RECT 92.390 50.690 92.665 50.750 ;
        RECT 97.725 50.690 98.000 50.750 ;
        RECT 103.050 50.690 103.325 50.750 ;
        RECT 108.385 50.690 108.660 50.750 ;
        RECT 113.710 50.690 113.985 50.750 ;
        RECT 119.045 50.690 119.320 50.750 ;
        RECT 32.195 49.880 32.455 50.575 ;
        RECT 35.335 49.785 35.595 50.575 ;
        RECT 122.800 50.575 124.040 50.805 ;
        RECT 124.315 50.750 124.705 51.170 ;
        RECT 124.960 51.115 126.200 51.345 ;
        RECT 124.370 50.690 124.645 50.750 ;
        RECT 124.960 50.575 126.200 50.805 ;
        RECT 122.800 49.880 123.060 50.575 ;
        RECT 125.940 49.785 126.200 50.575 ;
        RECT 32.195 43.810 32.455 44.690 ;
        RECT 35.335 43.810 35.595 44.600 ;
        RECT 32.195 43.580 33.435 43.810 ;
        RECT 33.765 43.635 34.040 43.700 ;
        RECT 32.195 43.040 33.435 43.270 ;
        RECT 33.710 43.215 34.100 43.635 ;
        RECT 34.355 43.580 35.595 43.810 ;
        RECT 122.800 43.810 123.060 44.690 ;
        RECT 125.940 43.810 126.200 44.600 ;
        RECT 39.090 43.635 39.365 43.700 ;
        RECT 44.425 43.635 44.700 43.700 ;
        RECT 49.750 43.635 50.025 43.700 ;
        RECT 55.085 43.635 55.360 43.700 ;
        RECT 60.410 43.635 60.685 43.700 ;
        RECT 65.745 43.635 66.020 43.700 ;
        RECT 71.070 43.635 71.345 43.700 ;
        RECT 76.405 43.635 76.680 43.700 ;
        RECT 81.730 43.635 82.005 43.700 ;
        RECT 87.065 43.635 87.340 43.700 ;
        RECT 92.390 43.635 92.665 43.700 ;
        RECT 97.725 43.635 98.000 43.700 ;
        RECT 103.050 43.635 103.325 43.700 ;
        RECT 108.385 43.635 108.660 43.700 ;
        RECT 113.710 43.635 113.985 43.700 ;
        RECT 119.045 43.635 119.320 43.700 ;
        RECT 33.765 43.155 34.040 43.215 ;
        RECT 34.355 43.040 35.595 43.270 ;
        RECT 39.035 43.215 39.425 43.635 ;
        RECT 44.370 43.215 44.760 43.635 ;
        RECT 49.695 43.215 50.085 43.635 ;
        RECT 55.030 43.215 55.420 43.635 ;
        RECT 60.355 43.215 60.745 43.635 ;
        RECT 65.690 43.215 66.080 43.635 ;
        RECT 71.015 43.215 71.405 43.635 ;
        RECT 76.350 43.215 76.740 43.635 ;
        RECT 81.675 43.215 82.065 43.635 ;
        RECT 87.010 43.215 87.400 43.635 ;
        RECT 92.335 43.215 92.725 43.635 ;
        RECT 97.670 43.215 98.060 43.635 ;
        RECT 102.995 43.215 103.385 43.635 ;
        RECT 108.330 43.215 108.720 43.635 ;
        RECT 113.655 43.215 114.045 43.635 ;
        RECT 118.990 43.215 119.380 43.635 ;
        RECT 122.800 43.580 124.040 43.810 ;
        RECT 124.370 43.635 124.645 43.700 ;
        RECT 39.090 43.155 39.365 43.215 ;
        RECT 44.425 43.155 44.700 43.215 ;
        RECT 49.750 43.155 50.025 43.215 ;
        RECT 55.085 43.155 55.360 43.215 ;
        RECT 60.410 43.155 60.685 43.215 ;
        RECT 65.745 43.155 66.020 43.215 ;
        RECT 71.070 43.155 71.345 43.215 ;
        RECT 76.405 43.155 76.680 43.215 ;
        RECT 81.730 43.155 82.005 43.215 ;
        RECT 87.065 43.155 87.340 43.215 ;
        RECT 92.390 43.155 92.665 43.215 ;
        RECT 97.725 43.155 98.000 43.215 ;
        RECT 103.050 43.155 103.325 43.215 ;
        RECT 108.385 43.155 108.660 43.215 ;
        RECT 113.710 43.155 113.985 43.215 ;
        RECT 119.045 43.155 119.320 43.215 ;
        RECT 32.195 42.345 32.455 43.040 ;
        RECT 35.335 42.250 35.595 43.040 ;
        RECT 122.800 43.040 124.040 43.270 ;
        RECT 124.315 43.215 124.705 43.635 ;
        RECT 124.960 43.580 126.200 43.810 ;
        RECT 124.370 43.155 124.645 43.215 ;
        RECT 124.960 43.040 126.200 43.270 ;
        RECT 122.800 42.345 123.060 43.040 ;
        RECT 125.940 42.250 126.200 43.040 ;
        RECT 32.195 36.275 32.455 37.155 ;
        RECT 35.335 36.275 35.595 37.065 ;
        RECT 32.195 36.045 33.435 36.275 ;
        RECT 33.765 36.100 34.040 36.165 ;
        RECT 32.195 35.505 33.435 35.735 ;
        RECT 33.710 35.680 34.100 36.100 ;
        RECT 34.355 36.045 35.595 36.275 ;
        RECT 122.800 36.275 123.060 37.155 ;
        RECT 125.940 36.275 126.200 37.065 ;
        RECT 39.090 36.100 39.365 36.165 ;
        RECT 44.425 36.100 44.700 36.165 ;
        RECT 49.750 36.100 50.025 36.165 ;
        RECT 55.085 36.100 55.360 36.165 ;
        RECT 60.410 36.100 60.685 36.165 ;
        RECT 65.745 36.100 66.020 36.165 ;
        RECT 71.070 36.100 71.345 36.165 ;
        RECT 76.405 36.100 76.680 36.165 ;
        RECT 81.730 36.100 82.005 36.165 ;
        RECT 87.065 36.100 87.340 36.165 ;
        RECT 92.390 36.100 92.665 36.165 ;
        RECT 97.725 36.100 98.000 36.165 ;
        RECT 103.050 36.100 103.325 36.165 ;
        RECT 108.385 36.100 108.660 36.165 ;
        RECT 113.710 36.100 113.985 36.165 ;
        RECT 119.045 36.100 119.320 36.165 ;
        RECT 33.765 35.620 34.040 35.680 ;
        RECT 34.355 35.505 35.595 35.735 ;
        RECT 39.035 35.680 39.425 36.100 ;
        RECT 44.370 35.680 44.760 36.100 ;
        RECT 49.695 35.680 50.085 36.100 ;
        RECT 55.030 35.680 55.420 36.100 ;
        RECT 60.355 35.680 60.745 36.100 ;
        RECT 65.690 35.680 66.080 36.100 ;
        RECT 71.015 35.680 71.405 36.100 ;
        RECT 76.350 35.680 76.740 36.100 ;
        RECT 81.675 35.680 82.065 36.100 ;
        RECT 87.010 35.680 87.400 36.100 ;
        RECT 92.335 35.680 92.725 36.100 ;
        RECT 97.670 35.680 98.060 36.100 ;
        RECT 102.995 35.680 103.385 36.100 ;
        RECT 108.330 35.680 108.720 36.100 ;
        RECT 113.655 35.680 114.045 36.100 ;
        RECT 118.990 35.680 119.380 36.100 ;
        RECT 122.800 36.045 124.040 36.275 ;
        RECT 124.370 36.100 124.645 36.165 ;
        RECT 39.090 35.620 39.365 35.680 ;
        RECT 44.425 35.620 44.700 35.680 ;
        RECT 49.750 35.620 50.025 35.680 ;
        RECT 55.085 35.620 55.360 35.680 ;
        RECT 60.410 35.620 60.685 35.680 ;
        RECT 65.745 35.620 66.020 35.680 ;
        RECT 71.070 35.620 71.345 35.680 ;
        RECT 76.405 35.620 76.680 35.680 ;
        RECT 81.730 35.620 82.005 35.680 ;
        RECT 87.065 35.620 87.340 35.680 ;
        RECT 92.390 35.620 92.665 35.680 ;
        RECT 97.725 35.620 98.000 35.680 ;
        RECT 103.050 35.620 103.325 35.680 ;
        RECT 108.385 35.620 108.660 35.680 ;
        RECT 113.710 35.620 113.985 35.680 ;
        RECT 119.045 35.620 119.320 35.680 ;
        RECT 32.195 34.810 32.455 35.505 ;
        RECT 35.335 34.715 35.595 35.505 ;
        RECT 122.800 35.505 124.040 35.735 ;
        RECT 124.315 35.680 124.705 36.100 ;
        RECT 124.960 36.045 126.200 36.275 ;
        RECT 124.370 35.620 124.645 35.680 ;
        RECT 124.960 35.505 126.200 35.735 ;
        RECT 122.800 34.810 123.060 35.505 ;
        RECT 125.940 34.715 126.200 35.505 ;
        RECT 32.195 28.740 32.455 29.620 ;
        RECT 35.335 28.740 35.595 29.530 ;
        RECT 32.195 28.510 33.435 28.740 ;
        RECT 33.765 28.565 34.040 28.630 ;
        RECT 32.195 27.970 33.435 28.200 ;
        RECT 33.710 28.145 34.100 28.565 ;
        RECT 34.355 28.510 35.595 28.740 ;
        RECT 122.800 28.740 123.060 29.620 ;
        RECT 125.940 28.740 126.200 29.530 ;
        RECT 39.090 28.565 39.365 28.630 ;
        RECT 44.425 28.565 44.700 28.630 ;
        RECT 49.750 28.565 50.025 28.630 ;
        RECT 55.085 28.565 55.360 28.630 ;
        RECT 60.410 28.565 60.685 28.630 ;
        RECT 65.745 28.565 66.020 28.630 ;
        RECT 71.070 28.565 71.345 28.630 ;
        RECT 76.405 28.565 76.680 28.630 ;
        RECT 81.730 28.565 82.005 28.630 ;
        RECT 87.065 28.565 87.340 28.630 ;
        RECT 92.390 28.565 92.665 28.630 ;
        RECT 97.725 28.565 98.000 28.630 ;
        RECT 103.050 28.565 103.325 28.630 ;
        RECT 108.385 28.565 108.660 28.630 ;
        RECT 113.710 28.565 113.985 28.630 ;
        RECT 119.045 28.565 119.320 28.630 ;
        RECT 33.765 28.085 34.040 28.145 ;
        RECT 34.355 27.970 35.595 28.200 ;
        RECT 39.035 28.145 39.425 28.565 ;
        RECT 44.370 28.145 44.760 28.565 ;
        RECT 49.695 28.145 50.085 28.565 ;
        RECT 55.030 28.145 55.420 28.565 ;
        RECT 60.355 28.145 60.745 28.565 ;
        RECT 65.690 28.145 66.080 28.565 ;
        RECT 71.015 28.145 71.405 28.565 ;
        RECT 76.350 28.145 76.740 28.565 ;
        RECT 81.675 28.145 82.065 28.565 ;
        RECT 87.010 28.145 87.400 28.565 ;
        RECT 92.335 28.145 92.725 28.565 ;
        RECT 97.670 28.145 98.060 28.565 ;
        RECT 102.995 28.145 103.385 28.565 ;
        RECT 108.330 28.145 108.720 28.565 ;
        RECT 113.655 28.145 114.045 28.565 ;
        RECT 118.990 28.145 119.380 28.565 ;
        RECT 122.800 28.510 124.040 28.740 ;
        RECT 124.370 28.565 124.645 28.630 ;
        RECT 39.090 28.085 39.365 28.145 ;
        RECT 44.425 28.085 44.700 28.145 ;
        RECT 49.750 28.085 50.025 28.145 ;
        RECT 55.085 28.085 55.360 28.145 ;
        RECT 60.410 28.085 60.685 28.145 ;
        RECT 65.745 28.085 66.020 28.145 ;
        RECT 71.070 28.085 71.345 28.145 ;
        RECT 76.405 28.085 76.680 28.145 ;
        RECT 81.730 28.085 82.005 28.145 ;
        RECT 87.065 28.085 87.340 28.145 ;
        RECT 92.390 28.085 92.665 28.145 ;
        RECT 97.725 28.085 98.000 28.145 ;
        RECT 103.050 28.085 103.325 28.145 ;
        RECT 108.385 28.085 108.660 28.145 ;
        RECT 113.710 28.085 113.985 28.145 ;
        RECT 119.045 28.085 119.320 28.145 ;
        RECT 32.195 27.275 32.455 27.970 ;
        RECT 35.335 27.180 35.595 27.970 ;
        RECT 122.800 27.970 124.040 28.200 ;
        RECT 124.315 28.145 124.705 28.565 ;
        RECT 124.960 28.510 126.200 28.740 ;
        RECT 124.370 28.085 124.645 28.145 ;
        RECT 124.960 27.970 126.200 28.200 ;
        RECT 122.800 27.275 123.060 27.970 ;
        RECT 125.940 27.180 126.200 27.970 ;
        RECT 32.195 21.205 32.455 22.085 ;
        RECT 35.335 21.205 35.595 21.995 ;
        RECT 32.195 20.975 33.435 21.205 ;
        RECT 33.765 21.030 34.040 21.095 ;
        RECT 32.195 20.435 33.435 20.665 ;
        RECT 33.710 20.610 34.100 21.030 ;
        RECT 34.355 20.975 35.595 21.205 ;
        RECT 122.800 21.205 123.060 22.085 ;
        RECT 125.940 21.205 126.200 21.995 ;
        RECT 39.090 21.030 39.365 21.095 ;
        RECT 44.425 21.030 44.700 21.095 ;
        RECT 49.750 21.030 50.025 21.095 ;
        RECT 55.085 21.030 55.360 21.095 ;
        RECT 60.410 21.030 60.685 21.095 ;
        RECT 65.745 21.030 66.020 21.095 ;
        RECT 71.070 21.030 71.345 21.095 ;
        RECT 76.405 21.030 76.680 21.095 ;
        RECT 81.730 21.030 82.005 21.095 ;
        RECT 87.065 21.030 87.340 21.095 ;
        RECT 92.390 21.030 92.665 21.095 ;
        RECT 97.725 21.030 98.000 21.095 ;
        RECT 103.050 21.030 103.325 21.095 ;
        RECT 108.385 21.030 108.660 21.095 ;
        RECT 113.710 21.030 113.985 21.095 ;
        RECT 119.045 21.030 119.320 21.095 ;
        RECT 33.765 20.550 34.040 20.610 ;
        RECT 34.355 20.435 35.595 20.665 ;
        RECT 39.035 20.610 39.425 21.030 ;
        RECT 44.370 20.610 44.760 21.030 ;
        RECT 49.695 20.610 50.085 21.030 ;
        RECT 55.030 20.610 55.420 21.030 ;
        RECT 60.355 20.610 60.745 21.030 ;
        RECT 65.690 20.610 66.080 21.030 ;
        RECT 71.015 20.610 71.405 21.030 ;
        RECT 76.350 20.610 76.740 21.030 ;
        RECT 81.675 20.610 82.065 21.030 ;
        RECT 87.010 20.610 87.400 21.030 ;
        RECT 92.335 20.610 92.725 21.030 ;
        RECT 97.670 20.610 98.060 21.030 ;
        RECT 102.995 20.610 103.385 21.030 ;
        RECT 108.330 20.610 108.720 21.030 ;
        RECT 113.655 20.610 114.045 21.030 ;
        RECT 118.990 20.610 119.380 21.030 ;
        RECT 122.800 20.975 124.040 21.205 ;
        RECT 124.370 21.030 124.645 21.095 ;
        RECT 39.090 20.550 39.365 20.610 ;
        RECT 44.425 20.550 44.700 20.610 ;
        RECT 49.750 20.550 50.025 20.610 ;
        RECT 55.085 20.550 55.360 20.610 ;
        RECT 60.410 20.550 60.685 20.610 ;
        RECT 65.745 20.550 66.020 20.610 ;
        RECT 71.070 20.550 71.345 20.610 ;
        RECT 76.405 20.550 76.680 20.610 ;
        RECT 81.730 20.550 82.005 20.610 ;
        RECT 87.065 20.550 87.340 20.610 ;
        RECT 92.390 20.550 92.665 20.610 ;
        RECT 97.725 20.550 98.000 20.610 ;
        RECT 103.050 20.550 103.325 20.610 ;
        RECT 108.385 20.550 108.660 20.610 ;
        RECT 113.710 20.550 113.985 20.610 ;
        RECT 119.045 20.550 119.320 20.610 ;
        RECT 32.195 19.740 32.455 20.435 ;
        RECT 35.335 19.645 35.595 20.435 ;
        RECT 122.800 20.435 124.040 20.665 ;
        RECT 124.315 20.610 124.705 21.030 ;
        RECT 124.960 20.975 126.200 21.205 ;
        RECT 124.370 20.550 124.645 20.610 ;
        RECT 124.960 20.435 126.200 20.665 ;
        RECT 122.800 19.740 123.060 20.435 ;
        RECT 125.940 19.645 126.200 20.435 ;
        RECT 32.195 13.670 32.455 14.550 ;
        RECT 35.335 13.670 35.595 14.460 ;
        RECT 32.195 13.440 33.435 13.670 ;
        RECT 33.765 13.495 34.040 13.560 ;
        RECT 32.195 12.900 33.435 13.130 ;
        RECT 33.710 13.075 34.100 13.495 ;
        RECT 34.355 13.440 35.595 13.670 ;
        RECT 122.800 13.670 123.060 14.550 ;
        RECT 125.940 13.670 126.200 14.460 ;
        RECT 39.090 13.495 39.365 13.560 ;
        RECT 44.425 13.495 44.700 13.560 ;
        RECT 49.750 13.495 50.025 13.560 ;
        RECT 55.085 13.495 55.360 13.560 ;
        RECT 60.410 13.495 60.685 13.560 ;
        RECT 65.745 13.495 66.020 13.560 ;
        RECT 71.070 13.495 71.345 13.560 ;
        RECT 76.405 13.495 76.680 13.560 ;
        RECT 81.730 13.495 82.005 13.560 ;
        RECT 87.065 13.495 87.340 13.560 ;
        RECT 92.390 13.495 92.665 13.560 ;
        RECT 97.725 13.495 98.000 13.560 ;
        RECT 103.050 13.495 103.325 13.560 ;
        RECT 108.385 13.495 108.660 13.560 ;
        RECT 113.710 13.495 113.985 13.560 ;
        RECT 119.045 13.495 119.320 13.560 ;
        RECT 33.765 13.015 34.040 13.075 ;
        RECT 34.355 12.900 35.595 13.130 ;
        RECT 39.035 13.075 39.425 13.495 ;
        RECT 44.370 13.075 44.760 13.495 ;
        RECT 49.695 13.075 50.085 13.495 ;
        RECT 55.030 13.075 55.420 13.495 ;
        RECT 60.355 13.075 60.745 13.495 ;
        RECT 65.690 13.075 66.080 13.495 ;
        RECT 71.015 13.075 71.405 13.495 ;
        RECT 76.350 13.075 76.740 13.495 ;
        RECT 81.675 13.075 82.065 13.495 ;
        RECT 87.010 13.075 87.400 13.495 ;
        RECT 92.335 13.075 92.725 13.495 ;
        RECT 97.670 13.075 98.060 13.495 ;
        RECT 102.995 13.075 103.385 13.495 ;
        RECT 108.330 13.075 108.720 13.495 ;
        RECT 113.655 13.075 114.045 13.495 ;
        RECT 118.990 13.075 119.380 13.495 ;
        RECT 122.800 13.440 124.040 13.670 ;
        RECT 124.370 13.495 124.645 13.560 ;
        RECT 39.090 13.015 39.365 13.075 ;
        RECT 44.425 13.015 44.700 13.075 ;
        RECT 49.750 13.015 50.025 13.075 ;
        RECT 55.085 13.015 55.360 13.075 ;
        RECT 60.410 13.015 60.685 13.075 ;
        RECT 65.745 13.015 66.020 13.075 ;
        RECT 71.070 13.015 71.345 13.075 ;
        RECT 76.405 13.015 76.680 13.075 ;
        RECT 81.730 13.015 82.005 13.075 ;
        RECT 87.065 13.015 87.340 13.075 ;
        RECT 92.390 13.015 92.665 13.075 ;
        RECT 97.725 13.015 98.000 13.075 ;
        RECT 103.050 13.015 103.325 13.075 ;
        RECT 108.385 13.015 108.660 13.075 ;
        RECT 113.710 13.015 113.985 13.075 ;
        RECT 119.045 13.015 119.320 13.075 ;
        RECT 32.195 12.205 32.455 12.900 ;
        RECT 35.335 12.110 35.595 12.900 ;
        RECT 122.800 12.900 124.040 13.130 ;
        RECT 124.315 13.075 124.705 13.495 ;
        RECT 124.960 13.440 126.200 13.670 ;
        RECT 124.370 13.015 124.645 13.075 ;
        RECT 124.960 12.900 126.200 13.130 ;
        RECT 122.800 12.205 123.060 12.900 ;
        RECT 125.940 12.110 126.200 12.900 ;
        RECT 32.195 6.135 32.455 7.015 ;
        RECT 35.335 6.135 35.595 6.925 ;
        RECT 32.195 5.905 33.435 6.135 ;
        RECT 33.765 5.960 34.040 6.025 ;
        RECT 32.195 5.365 33.435 5.595 ;
        RECT 33.710 5.540 34.100 5.960 ;
        RECT 34.355 5.905 35.595 6.135 ;
        RECT 37.520 6.135 37.780 7.015 ;
        RECT 40.660 6.135 40.920 6.925 ;
        RECT 37.520 5.905 38.760 6.135 ;
        RECT 39.090 5.960 39.365 6.025 ;
        RECT 33.765 5.480 34.040 5.540 ;
        RECT 34.355 5.365 35.595 5.595 ;
        RECT 32.195 4.670 32.455 5.365 ;
        RECT 35.335 4.575 35.595 5.365 ;
        RECT 37.520 5.365 38.760 5.595 ;
        RECT 39.035 5.540 39.425 5.960 ;
        RECT 39.680 5.905 40.920 6.135 ;
        RECT 42.855 6.135 43.115 7.015 ;
        RECT 45.995 6.135 46.255 6.925 ;
        RECT 42.855 5.905 44.095 6.135 ;
        RECT 44.425 5.960 44.700 6.025 ;
        RECT 39.090 5.480 39.365 5.540 ;
        RECT 39.680 5.365 40.920 5.595 ;
        RECT 37.520 4.670 37.780 5.365 ;
        RECT 40.660 4.575 40.920 5.365 ;
        RECT 42.855 5.365 44.095 5.595 ;
        RECT 44.370 5.540 44.760 5.960 ;
        RECT 45.015 5.905 46.255 6.135 ;
        RECT 48.180 6.135 48.440 7.015 ;
        RECT 51.320 6.135 51.580 6.925 ;
        RECT 48.180 5.905 49.420 6.135 ;
        RECT 49.750 5.960 50.025 6.025 ;
        RECT 44.425 5.480 44.700 5.540 ;
        RECT 45.015 5.365 46.255 5.595 ;
        RECT 42.855 4.670 43.115 5.365 ;
        RECT 45.995 4.575 46.255 5.365 ;
        RECT 48.180 5.365 49.420 5.595 ;
        RECT 49.695 5.540 50.085 5.960 ;
        RECT 50.340 5.905 51.580 6.135 ;
        RECT 53.515 6.135 53.775 7.015 ;
        RECT 56.655 6.135 56.915 6.925 ;
        RECT 53.515 5.905 54.755 6.135 ;
        RECT 55.085 5.960 55.360 6.025 ;
        RECT 49.750 5.480 50.025 5.540 ;
        RECT 50.340 5.365 51.580 5.595 ;
        RECT 48.180 4.670 48.440 5.365 ;
        RECT 51.320 4.575 51.580 5.365 ;
        RECT 53.515 5.365 54.755 5.595 ;
        RECT 55.030 5.540 55.420 5.960 ;
        RECT 55.675 5.905 56.915 6.135 ;
        RECT 58.840 6.135 59.100 7.015 ;
        RECT 61.980 6.135 62.240 6.925 ;
        RECT 58.840 5.905 60.080 6.135 ;
        RECT 60.410 5.960 60.685 6.025 ;
        RECT 55.085 5.480 55.360 5.540 ;
        RECT 55.675 5.365 56.915 5.595 ;
        RECT 53.515 4.670 53.775 5.365 ;
        RECT 56.655 4.575 56.915 5.365 ;
        RECT 58.840 5.365 60.080 5.595 ;
        RECT 60.355 5.540 60.745 5.960 ;
        RECT 61.000 5.905 62.240 6.135 ;
        RECT 64.175 6.135 64.435 7.015 ;
        RECT 67.315 6.135 67.575 6.925 ;
        RECT 64.175 5.905 65.415 6.135 ;
        RECT 65.745 5.960 66.020 6.025 ;
        RECT 60.410 5.480 60.685 5.540 ;
        RECT 61.000 5.365 62.240 5.595 ;
        RECT 58.840 4.670 59.100 5.365 ;
        RECT 61.980 4.575 62.240 5.365 ;
        RECT 64.175 5.365 65.415 5.595 ;
        RECT 65.690 5.540 66.080 5.960 ;
        RECT 66.335 5.905 67.575 6.135 ;
        RECT 69.500 6.135 69.760 7.015 ;
        RECT 72.640 6.135 72.900 6.925 ;
        RECT 69.500 5.905 70.740 6.135 ;
        RECT 71.070 5.960 71.345 6.025 ;
        RECT 65.745 5.480 66.020 5.540 ;
        RECT 66.335 5.365 67.575 5.595 ;
        RECT 64.175 4.670 64.435 5.365 ;
        RECT 67.315 4.575 67.575 5.365 ;
        RECT 69.500 5.365 70.740 5.595 ;
        RECT 71.015 5.540 71.405 5.960 ;
        RECT 71.660 5.905 72.900 6.135 ;
        RECT 74.835 6.135 75.095 7.015 ;
        RECT 77.975 6.135 78.235 6.925 ;
        RECT 74.835 5.905 76.075 6.135 ;
        RECT 76.405 5.960 76.680 6.025 ;
        RECT 71.070 5.480 71.345 5.540 ;
        RECT 71.660 5.365 72.900 5.595 ;
        RECT 69.500 4.670 69.760 5.365 ;
        RECT 72.640 4.575 72.900 5.365 ;
        RECT 74.835 5.365 76.075 5.595 ;
        RECT 76.350 5.540 76.740 5.960 ;
        RECT 76.995 5.905 78.235 6.135 ;
        RECT 80.160 6.135 80.420 7.015 ;
        RECT 83.300 6.135 83.560 6.925 ;
        RECT 80.160 5.905 81.400 6.135 ;
        RECT 81.730 5.960 82.005 6.025 ;
        RECT 76.405 5.480 76.680 5.540 ;
        RECT 76.995 5.365 78.235 5.595 ;
        RECT 74.835 4.670 75.095 5.365 ;
        RECT 77.975 4.575 78.235 5.365 ;
        RECT 80.160 5.365 81.400 5.595 ;
        RECT 81.675 5.540 82.065 5.960 ;
        RECT 82.320 5.905 83.560 6.135 ;
        RECT 85.495 6.135 85.755 7.015 ;
        RECT 88.635 6.135 88.895 6.925 ;
        RECT 85.495 5.905 86.735 6.135 ;
        RECT 87.065 5.960 87.340 6.025 ;
        RECT 81.730 5.480 82.005 5.540 ;
        RECT 82.320 5.365 83.560 5.595 ;
        RECT 80.160 4.670 80.420 5.365 ;
        RECT 83.300 4.575 83.560 5.365 ;
        RECT 85.495 5.365 86.735 5.595 ;
        RECT 87.010 5.540 87.400 5.960 ;
        RECT 87.655 5.905 88.895 6.135 ;
        RECT 90.820 6.135 91.080 7.015 ;
        RECT 93.960 6.135 94.220 6.925 ;
        RECT 90.820 5.905 92.060 6.135 ;
        RECT 92.390 5.960 92.665 6.025 ;
        RECT 87.065 5.480 87.340 5.540 ;
        RECT 87.655 5.365 88.895 5.595 ;
        RECT 85.495 4.670 85.755 5.365 ;
        RECT 88.635 4.575 88.895 5.365 ;
        RECT 90.820 5.365 92.060 5.595 ;
        RECT 92.335 5.540 92.725 5.960 ;
        RECT 92.980 5.905 94.220 6.135 ;
        RECT 96.155 6.135 96.415 7.015 ;
        RECT 99.295 6.135 99.555 6.925 ;
        RECT 96.155 5.905 97.395 6.135 ;
        RECT 97.725 5.960 98.000 6.025 ;
        RECT 92.390 5.480 92.665 5.540 ;
        RECT 92.980 5.365 94.220 5.595 ;
        RECT 90.820 4.670 91.080 5.365 ;
        RECT 93.960 4.575 94.220 5.365 ;
        RECT 96.155 5.365 97.395 5.595 ;
        RECT 97.670 5.540 98.060 5.960 ;
        RECT 98.315 5.905 99.555 6.135 ;
        RECT 101.480 6.135 101.740 7.015 ;
        RECT 104.620 6.135 104.880 6.925 ;
        RECT 101.480 5.905 102.720 6.135 ;
        RECT 103.050 5.960 103.325 6.025 ;
        RECT 97.725 5.480 98.000 5.540 ;
        RECT 98.315 5.365 99.555 5.595 ;
        RECT 96.155 4.670 96.415 5.365 ;
        RECT 99.295 4.575 99.555 5.365 ;
        RECT 101.480 5.365 102.720 5.595 ;
        RECT 102.995 5.540 103.385 5.960 ;
        RECT 103.640 5.905 104.880 6.135 ;
        RECT 106.815 6.135 107.075 7.015 ;
        RECT 109.955 6.135 110.215 6.925 ;
        RECT 106.815 5.905 108.055 6.135 ;
        RECT 108.385 5.960 108.660 6.025 ;
        RECT 103.050 5.480 103.325 5.540 ;
        RECT 103.640 5.365 104.880 5.595 ;
        RECT 101.480 4.670 101.740 5.365 ;
        RECT 104.620 4.575 104.880 5.365 ;
        RECT 106.815 5.365 108.055 5.595 ;
        RECT 108.330 5.540 108.720 5.960 ;
        RECT 108.975 5.905 110.215 6.135 ;
        RECT 112.140 6.135 112.400 7.015 ;
        RECT 115.280 6.135 115.540 6.925 ;
        RECT 112.140 5.905 113.380 6.135 ;
        RECT 113.710 5.960 113.985 6.025 ;
        RECT 108.385 5.480 108.660 5.540 ;
        RECT 108.975 5.365 110.215 5.595 ;
        RECT 106.815 4.670 107.075 5.365 ;
        RECT 109.955 4.575 110.215 5.365 ;
        RECT 112.140 5.365 113.380 5.595 ;
        RECT 113.655 5.540 114.045 5.960 ;
        RECT 114.300 5.905 115.540 6.135 ;
        RECT 117.475 6.135 117.735 7.015 ;
        RECT 120.615 6.135 120.875 6.925 ;
        RECT 117.475 5.905 118.715 6.135 ;
        RECT 119.045 5.960 119.320 6.025 ;
        RECT 113.710 5.480 113.985 5.540 ;
        RECT 114.300 5.365 115.540 5.595 ;
        RECT 112.140 4.670 112.400 5.365 ;
        RECT 115.280 4.575 115.540 5.365 ;
        RECT 117.475 5.365 118.715 5.595 ;
        RECT 118.990 5.540 119.380 5.960 ;
        RECT 119.635 5.905 120.875 6.135 ;
        RECT 122.800 6.135 123.060 7.015 ;
        RECT 125.940 6.135 126.200 6.925 ;
        RECT 122.800 5.905 124.040 6.135 ;
        RECT 124.370 5.960 124.645 6.025 ;
        RECT 119.045 5.480 119.320 5.540 ;
        RECT 119.635 5.365 120.875 5.595 ;
        RECT 117.475 4.670 117.735 5.365 ;
        RECT 120.615 4.575 120.875 5.365 ;
        RECT 122.800 5.365 124.040 5.595 ;
        RECT 124.315 5.540 124.705 5.960 ;
        RECT 124.960 5.905 126.200 6.135 ;
        RECT 124.370 5.480 124.645 5.540 ;
        RECT 124.960 5.365 126.200 5.595 ;
        RECT 122.800 4.670 123.060 5.365 ;
        RECT 125.940 4.575 126.200 5.365 ;
      LAYER met2 ;
        RECT 62.035 84.500 63.845 84.510 ;
        RECT 66.480 84.500 68.385 84.510 ;
        RECT 71.025 84.500 74.615 84.510 ;
        RECT 62.035 81.815 74.615 84.500 ;
        RECT 29.785 74.155 30.925 78.295 ;
        RECT 31.460 74.800 31.830 74.810 ;
        RECT 36.785 74.800 37.155 74.810 ;
        RECT 42.120 74.800 42.490 74.810 ;
        RECT 47.445 74.800 47.815 74.810 ;
        RECT 52.780 74.800 53.150 74.810 ;
        RECT 58.105 74.800 58.475 74.810 ;
        RECT 63.440 74.800 63.810 74.810 ;
        RECT 68.765 74.800 69.135 74.810 ;
        RECT 74.100 74.800 74.470 74.810 ;
        RECT 79.425 74.800 79.795 74.810 ;
        RECT 84.760 74.800 85.130 74.810 ;
        RECT 90.085 74.800 90.455 74.810 ;
        RECT 95.420 74.800 95.790 74.810 ;
        RECT 100.745 74.800 101.115 74.810 ;
        RECT 106.080 74.800 106.450 74.810 ;
        RECT 111.405 74.800 111.775 74.810 ;
        RECT 116.740 74.800 117.110 74.810 ;
        RECT 122.065 74.800 122.435 74.810 ;
        RECT 31.460 74.540 32.485 74.800 ;
        RECT 35.960 74.710 36.330 74.720 ;
        RECT 31.460 74.530 31.830 74.540 ;
        RECT 32.195 74.155 32.455 74.540 ;
        RECT 35.305 74.450 36.330 74.710 ;
        RECT 36.785 74.540 37.810 74.800 ;
        RECT 41.285 74.710 41.655 74.720 ;
        RECT 36.785 74.530 37.155 74.540 ;
        RECT 35.335 74.155 35.595 74.450 ;
        RECT 35.960 74.440 36.330 74.450 ;
        RECT 37.520 74.155 37.780 74.540 ;
        RECT 40.630 74.450 41.655 74.710 ;
        RECT 42.120 74.540 43.145 74.800 ;
        RECT 46.620 74.710 46.990 74.720 ;
        RECT 42.120 74.530 42.490 74.540 ;
        RECT 40.660 74.155 40.920 74.450 ;
        RECT 41.285 74.440 41.655 74.450 ;
        RECT 42.855 74.155 43.115 74.540 ;
        RECT 45.965 74.450 46.990 74.710 ;
        RECT 47.445 74.540 48.470 74.800 ;
        RECT 51.945 74.710 52.315 74.720 ;
        RECT 47.445 74.530 47.815 74.540 ;
        RECT 45.995 74.155 46.255 74.450 ;
        RECT 46.620 74.440 46.990 74.450 ;
        RECT 48.180 74.155 48.440 74.540 ;
        RECT 51.290 74.450 52.315 74.710 ;
        RECT 52.780 74.540 53.805 74.800 ;
        RECT 57.280 74.710 57.650 74.720 ;
        RECT 52.780 74.530 53.150 74.540 ;
        RECT 51.320 74.155 51.580 74.450 ;
        RECT 51.945 74.440 52.315 74.450 ;
        RECT 53.515 74.155 53.775 74.540 ;
        RECT 56.625 74.450 57.650 74.710 ;
        RECT 58.105 74.540 59.130 74.800 ;
        RECT 62.605 74.710 62.975 74.720 ;
        RECT 58.105 74.530 58.475 74.540 ;
        RECT 56.655 74.155 56.915 74.450 ;
        RECT 57.280 74.440 57.650 74.450 ;
        RECT 58.840 74.155 59.100 74.540 ;
        RECT 61.950 74.450 62.975 74.710 ;
        RECT 63.440 74.540 64.465 74.800 ;
        RECT 67.940 74.710 68.310 74.720 ;
        RECT 63.440 74.530 63.810 74.540 ;
        RECT 61.980 74.155 62.240 74.450 ;
        RECT 62.605 74.440 62.975 74.450 ;
        RECT 64.175 74.155 64.435 74.540 ;
        RECT 67.285 74.450 68.310 74.710 ;
        RECT 68.765 74.540 69.790 74.800 ;
        RECT 73.265 74.710 73.635 74.720 ;
        RECT 68.765 74.530 69.135 74.540 ;
        RECT 67.315 74.155 67.575 74.450 ;
        RECT 67.940 74.440 68.310 74.450 ;
        RECT 69.500 74.155 69.760 74.540 ;
        RECT 72.610 74.450 73.635 74.710 ;
        RECT 74.100 74.540 75.125 74.800 ;
        RECT 78.600 74.710 78.970 74.720 ;
        RECT 74.100 74.530 74.470 74.540 ;
        RECT 72.640 74.155 72.900 74.450 ;
        RECT 73.265 74.440 73.635 74.450 ;
        RECT 74.835 74.155 75.095 74.540 ;
        RECT 77.945 74.450 78.970 74.710 ;
        RECT 79.425 74.540 80.450 74.800 ;
        RECT 83.925 74.710 84.295 74.720 ;
        RECT 79.425 74.530 79.795 74.540 ;
        RECT 77.975 74.155 78.235 74.450 ;
        RECT 78.600 74.440 78.970 74.450 ;
        RECT 80.160 74.155 80.420 74.540 ;
        RECT 83.270 74.450 84.295 74.710 ;
        RECT 84.760 74.540 85.785 74.800 ;
        RECT 89.260 74.710 89.630 74.720 ;
        RECT 84.760 74.530 85.130 74.540 ;
        RECT 83.300 74.155 83.560 74.450 ;
        RECT 83.925 74.440 84.295 74.450 ;
        RECT 85.495 74.155 85.755 74.540 ;
        RECT 88.605 74.450 89.630 74.710 ;
        RECT 90.085 74.540 91.110 74.800 ;
        RECT 94.585 74.710 94.955 74.720 ;
        RECT 90.085 74.530 90.455 74.540 ;
        RECT 88.635 74.155 88.895 74.450 ;
        RECT 89.260 74.440 89.630 74.450 ;
        RECT 90.820 74.155 91.080 74.540 ;
        RECT 93.930 74.450 94.955 74.710 ;
        RECT 95.420 74.540 96.445 74.800 ;
        RECT 99.920 74.710 100.290 74.720 ;
        RECT 95.420 74.530 95.790 74.540 ;
        RECT 93.960 74.155 94.220 74.450 ;
        RECT 94.585 74.440 94.955 74.450 ;
        RECT 96.155 74.155 96.415 74.540 ;
        RECT 99.265 74.450 100.290 74.710 ;
        RECT 100.745 74.540 101.770 74.800 ;
        RECT 105.245 74.710 105.615 74.720 ;
        RECT 100.745 74.530 101.115 74.540 ;
        RECT 99.295 74.155 99.555 74.450 ;
        RECT 99.920 74.440 100.290 74.450 ;
        RECT 101.480 74.155 101.740 74.540 ;
        RECT 104.590 74.450 105.615 74.710 ;
        RECT 106.080 74.540 107.105 74.800 ;
        RECT 110.580 74.710 110.950 74.720 ;
        RECT 106.080 74.530 106.450 74.540 ;
        RECT 104.620 74.155 104.880 74.450 ;
        RECT 105.245 74.440 105.615 74.450 ;
        RECT 106.815 74.155 107.075 74.540 ;
        RECT 109.925 74.450 110.950 74.710 ;
        RECT 111.405 74.540 112.430 74.800 ;
        RECT 115.905 74.710 116.275 74.720 ;
        RECT 111.405 74.530 111.775 74.540 ;
        RECT 109.955 74.155 110.215 74.450 ;
        RECT 110.580 74.440 110.950 74.450 ;
        RECT 112.140 74.155 112.400 74.540 ;
        RECT 115.250 74.450 116.275 74.710 ;
        RECT 116.740 74.540 117.765 74.800 ;
        RECT 121.240 74.710 121.610 74.720 ;
        RECT 116.740 74.530 117.110 74.540 ;
        RECT 115.280 74.155 115.540 74.450 ;
        RECT 115.905 74.440 116.275 74.450 ;
        RECT 117.475 74.155 117.735 74.540 ;
        RECT 120.585 74.450 121.610 74.710 ;
        RECT 122.065 74.540 123.090 74.800 ;
        RECT 126.565 74.710 126.935 74.720 ;
        RECT 122.065 74.530 122.435 74.540 ;
        RECT 120.615 74.155 120.875 74.450 ;
        RECT 121.240 74.440 121.610 74.450 ;
        RECT 122.800 74.155 123.060 74.540 ;
        RECT 125.910 74.450 126.935 74.710 ;
        RECT 125.940 74.155 126.200 74.450 ;
        RECT 126.565 74.440 126.935 74.450 ;
        RECT 29.785 73.030 127.180 74.155 ;
        RECT 29.785 66.620 30.925 73.030 ;
        RECT 31.460 72.775 31.830 72.785 ;
        RECT 32.195 72.775 32.455 73.030 ;
        RECT 31.460 72.515 32.485 72.775 ;
        RECT 35.335 72.680 35.595 73.030 ;
        RECT 36.785 72.775 37.155 72.785 ;
        RECT 37.520 72.775 37.780 73.030 ;
        RECT 35.960 72.680 36.330 72.690 ;
        RECT 31.460 72.505 31.830 72.515 ;
        RECT 35.305 72.420 36.330 72.680 ;
        RECT 36.785 72.515 37.810 72.775 ;
        RECT 40.660 72.680 40.920 73.030 ;
        RECT 42.120 72.775 42.490 72.785 ;
        RECT 42.855 72.775 43.140 73.030 ;
        RECT 41.285 72.680 41.655 72.690 ;
        RECT 36.785 72.505 37.155 72.515 ;
        RECT 40.630 72.420 41.655 72.680 ;
        RECT 42.120 72.515 43.145 72.775 ;
        RECT 45.995 72.680 46.255 73.030 ;
        RECT 47.445 72.775 47.815 72.785 ;
        RECT 48.180 72.775 48.440 73.030 ;
        RECT 46.620 72.680 46.990 72.690 ;
        RECT 42.120 72.505 42.490 72.515 ;
        RECT 45.965 72.420 46.990 72.680 ;
        RECT 47.445 72.515 48.470 72.775 ;
        RECT 51.320 72.680 51.580 73.030 ;
        RECT 52.780 72.775 53.150 72.785 ;
        RECT 53.515 72.775 53.800 73.030 ;
        RECT 51.945 72.680 52.315 72.690 ;
        RECT 47.445 72.505 47.815 72.515 ;
        RECT 51.290 72.420 52.315 72.680 ;
        RECT 52.780 72.515 53.805 72.775 ;
        RECT 56.655 72.680 56.915 73.030 ;
        RECT 58.105 72.775 58.475 72.785 ;
        RECT 58.840 72.775 59.100 73.030 ;
        RECT 57.280 72.680 57.650 72.690 ;
        RECT 52.780 72.505 53.150 72.515 ;
        RECT 56.625 72.420 57.650 72.680 ;
        RECT 58.105 72.515 59.130 72.775 ;
        RECT 61.980 72.680 62.240 73.030 ;
        RECT 63.440 72.775 63.810 72.785 ;
        RECT 64.175 72.775 64.460 73.030 ;
        RECT 62.605 72.680 62.975 72.690 ;
        RECT 58.105 72.505 58.475 72.515 ;
        RECT 61.950 72.420 62.975 72.680 ;
        RECT 63.440 72.515 64.465 72.775 ;
        RECT 67.315 72.680 67.575 73.030 ;
        RECT 68.765 72.775 69.135 72.785 ;
        RECT 69.500 72.775 69.760 73.030 ;
        RECT 67.940 72.680 68.310 72.690 ;
        RECT 63.440 72.505 63.810 72.515 ;
        RECT 67.285 72.420 68.310 72.680 ;
        RECT 68.765 72.515 69.790 72.775 ;
        RECT 72.640 72.680 72.900 73.030 ;
        RECT 74.100 72.775 74.470 72.785 ;
        RECT 74.835 72.775 75.120 73.030 ;
        RECT 73.265 72.680 73.635 72.690 ;
        RECT 68.765 72.505 69.135 72.515 ;
        RECT 72.610 72.420 73.635 72.680 ;
        RECT 74.100 72.515 75.125 72.775 ;
        RECT 77.975 72.680 78.235 73.030 ;
        RECT 79.425 72.775 79.795 72.785 ;
        RECT 80.160 72.775 80.420 73.030 ;
        RECT 78.600 72.680 78.970 72.690 ;
        RECT 74.100 72.505 74.470 72.515 ;
        RECT 77.945 72.420 78.970 72.680 ;
        RECT 79.425 72.515 80.450 72.775 ;
        RECT 83.300 72.680 83.560 73.030 ;
        RECT 84.760 72.775 85.130 72.785 ;
        RECT 85.495 72.775 85.780 73.030 ;
        RECT 83.925 72.680 84.295 72.690 ;
        RECT 79.425 72.505 79.795 72.515 ;
        RECT 83.270 72.420 84.295 72.680 ;
        RECT 84.760 72.515 85.785 72.775 ;
        RECT 88.635 72.680 88.895 73.030 ;
        RECT 90.085 72.775 90.455 72.785 ;
        RECT 90.820 72.775 91.080 73.030 ;
        RECT 89.260 72.680 89.630 72.690 ;
        RECT 84.760 72.505 85.130 72.515 ;
        RECT 88.605 72.420 89.630 72.680 ;
        RECT 90.085 72.515 91.110 72.775 ;
        RECT 93.960 72.680 94.220 73.030 ;
        RECT 95.420 72.775 95.790 72.785 ;
        RECT 96.155 72.775 96.440 73.030 ;
        RECT 94.585 72.680 94.955 72.690 ;
        RECT 90.085 72.505 90.455 72.515 ;
        RECT 93.930 72.420 94.955 72.680 ;
        RECT 95.420 72.515 96.445 72.775 ;
        RECT 99.295 72.680 99.555 73.030 ;
        RECT 100.745 72.775 101.115 72.785 ;
        RECT 101.480 72.775 101.740 73.030 ;
        RECT 99.920 72.680 100.290 72.690 ;
        RECT 95.420 72.505 95.790 72.515 ;
        RECT 99.265 72.420 100.290 72.680 ;
        RECT 100.745 72.515 101.770 72.775 ;
        RECT 104.620 72.680 104.880 73.030 ;
        RECT 106.080 72.775 106.450 72.785 ;
        RECT 106.815 72.775 107.100 73.030 ;
        RECT 105.245 72.680 105.615 72.690 ;
        RECT 100.745 72.505 101.115 72.515 ;
        RECT 104.590 72.420 105.615 72.680 ;
        RECT 106.080 72.515 107.105 72.775 ;
        RECT 109.955 72.680 110.215 73.030 ;
        RECT 111.405 72.775 111.775 72.785 ;
        RECT 112.140 72.775 112.400 73.030 ;
        RECT 110.580 72.680 110.950 72.690 ;
        RECT 106.080 72.505 106.450 72.515 ;
        RECT 109.925 72.420 110.950 72.680 ;
        RECT 111.405 72.515 112.430 72.775 ;
        RECT 115.280 72.680 115.540 73.030 ;
        RECT 116.740 72.775 117.110 72.785 ;
        RECT 117.475 72.775 117.760 73.030 ;
        RECT 115.905 72.680 116.275 72.690 ;
        RECT 111.405 72.505 111.775 72.515 ;
        RECT 115.250 72.420 116.275 72.680 ;
        RECT 116.740 72.515 117.765 72.775 ;
        RECT 120.615 72.680 120.875 73.030 ;
        RECT 122.065 72.775 122.435 72.785 ;
        RECT 122.800 72.775 123.060 73.030 ;
        RECT 121.240 72.680 121.610 72.690 ;
        RECT 116.740 72.505 117.110 72.515 ;
        RECT 120.585 72.420 121.610 72.680 ;
        RECT 122.065 72.515 123.090 72.775 ;
        RECT 125.940 72.680 126.200 73.030 ;
        RECT 126.565 72.680 126.935 72.690 ;
        RECT 122.065 72.505 122.435 72.515 ;
        RECT 125.910 72.420 126.935 72.680 ;
        RECT 35.960 72.410 36.330 72.420 ;
        RECT 41.285 72.410 41.655 72.420 ;
        RECT 46.620 72.410 46.990 72.420 ;
        RECT 51.945 72.410 52.315 72.420 ;
        RECT 57.280 72.410 57.650 72.420 ;
        RECT 62.605 72.410 62.975 72.420 ;
        RECT 67.940 72.410 68.310 72.420 ;
        RECT 73.265 72.410 73.635 72.420 ;
        RECT 78.600 72.410 78.970 72.420 ;
        RECT 83.925 72.410 84.295 72.420 ;
        RECT 89.260 72.410 89.630 72.420 ;
        RECT 94.585 72.410 94.955 72.420 ;
        RECT 99.920 72.410 100.290 72.420 ;
        RECT 105.245 72.410 105.615 72.420 ;
        RECT 110.580 72.410 110.950 72.420 ;
        RECT 115.905 72.410 116.275 72.420 ;
        RECT 121.240 72.410 121.610 72.420 ;
        RECT 126.565 72.410 126.935 72.420 ;
        RECT 31.460 67.265 31.830 67.275 ;
        RECT 74.100 67.265 74.470 67.275 ;
        RECT 116.740 67.265 117.110 67.275 ;
        RECT 122.065 67.265 122.435 67.275 ;
        RECT 31.460 67.005 32.485 67.265 ;
        RECT 35.960 67.175 36.330 67.185 ;
        RECT 31.460 66.995 31.830 67.005 ;
        RECT 32.195 66.620 32.455 67.005 ;
        RECT 35.305 66.915 36.330 67.175 ;
        RECT 74.100 67.005 75.125 67.265 ;
        RECT 116.740 67.005 117.765 67.265 ;
        RECT 122.065 67.005 123.090 67.265 ;
        RECT 126.565 67.175 126.935 67.185 ;
        RECT 74.100 66.995 74.470 67.005 ;
        RECT 116.740 66.995 117.110 67.005 ;
        RECT 122.065 66.995 122.435 67.005 ;
        RECT 35.335 66.620 35.595 66.915 ;
        RECT 35.960 66.905 36.330 66.915 ;
        RECT 122.800 66.620 123.060 67.005 ;
        RECT 125.910 66.915 126.935 67.175 ;
        RECT 125.940 66.620 126.200 66.915 ;
        RECT 126.565 66.905 126.935 66.915 ;
        RECT 29.785 65.495 127.180 66.620 ;
        RECT 29.785 59.085 30.925 65.495 ;
        RECT 31.460 65.240 31.830 65.250 ;
        RECT 32.195 65.240 32.455 65.495 ;
        RECT 31.460 64.980 32.485 65.240 ;
        RECT 35.335 65.145 35.595 65.495 ;
        RECT 122.065 65.240 122.435 65.250 ;
        RECT 122.800 65.240 123.060 65.495 ;
        RECT 35.960 65.145 36.330 65.155 ;
        RECT 31.460 64.970 31.830 64.980 ;
        RECT 35.305 64.885 36.330 65.145 ;
        RECT 122.065 64.980 123.090 65.240 ;
        RECT 125.940 65.145 126.200 65.495 ;
        RECT 126.565 65.145 126.935 65.155 ;
        RECT 122.065 64.970 122.435 64.980 ;
        RECT 125.910 64.885 126.935 65.145 ;
        RECT 35.960 64.875 36.330 64.885 ;
        RECT 126.565 64.875 126.935 64.885 ;
        RECT 31.460 59.730 31.830 59.740 ;
        RECT 122.065 59.730 122.435 59.740 ;
        RECT 31.460 59.470 32.485 59.730 ;
        RECT 35.960 59.640 36.330 59.650 ;
        RECT 31.460 59.460 31.830 59.470 ;
        RECT 32.195 59.085 32.455 59.470 ;
        RECT 35.305 59.380 36.330 59.640 ;
        RECT 122.065 59.470 123.090 59.730 ;
        RECT 126.565 59.640 126.935 59.650 ;
        RECT 122.065 59.460 122.435 59.470 ;
        RECT 35.335 59.085 35.595 59.380 ;
        RECT 35.960 59.370 36.330 59.380 ;
        RECT 122.800 59.085 123.060 59.470 ;
        RECT 125.910 59.380 126.935 59.640 ;
        RECT 125.940 59.085 126.200 59.380 ;
        RECT 126.565 59.370 126.935 59.380 ;
        RECT 29.785 57.960 127.180 59.085 ;
        RECT 29.785 51.550 30.925 57.960 ;
        RECT 31.460 57.705 31.830 57.715 ;
        RECT 32.195 57.705 32.455 57.960 ;
        RECT 31.460 57.445 32.485 57.705 ;
        RECT 35.335 57.610 35.595 57.960 ;
        RECT 122.065 57.705 122.435 57.715 ;
        RECT 122.800 57.705 123.060 57.960 ;
        RECT 35.960 57.610 36.330 57.620 ;
        RECT 31.460 57.435 31.830 57.445 ;
        RECT 35.305 57.350 36.330 57.610 ;
        RECT 122.065 57.445 123.090 57.705 ;
        RECT 125.940 57.610 126.200 57.960 ;
        RECT 126.565 57.610 126.935 57.620 ;
        RECT 122.065 57.435 122.435 57.445 ;
        RECT 125.910 57.350 126.935 57.610 ;
        RECT 35.960 57.340 36.330 57.350 ;
        RECT 126.565 57.340 126.935 57.350 ;
        RECT 31.460 52.195 31.830 52.205 ;
        RECT 122.065 52.195 122.435 52.205 ;
        RECT 31.460 51.935 32.485 52.195 ;
        RECT 35.960 52.105 36.330 52.115 ;
        RECT 31.460 51.925 31.830 51.935 ;
        RECT 32.195 51.550 32.455 51.935 ;
        RECT 35.305 51.845 36.330 52.105 ;
        RECT 122.065 51.935 123.090 52.195 ;
        RECT 126.565 52.105 126.935 52.115 ;
        RECT 122.065 51.925 122.435 51.935 ;
        RECT 35.335 51.550 35.595 51.845 ;
        RECT 35.960 51.835 36.330 51.845 ;
        RECT 122.800 51.550 123.060 51.935 ;
        RECT 125.910 51.845 126.935 52.105 ;
        RECT 125.940 51.550 126.200 51.845 ;
        RECT 126.565 51.835 126.935 51.845 ;
        RECT 29.785 50.425 127.180 51.550 ;
        RECT 29.785 44.015 30.925 50.425 ;
        RECT 31.460 50.170 31.830 50.180 ;
        RECT 32.195 50.170 32.455 50.425 ;
        RECT 31.460 49.910 32.485 50.170 ;
        RECT 35.335 50.075 35.595 50.425 ;
        RECT 122.065 50.170 122.435 50.180 ;
        RECT 122.800 50.170 123.060 50.425 ;
        RECT 35.960 50.075 36.330 50.085 ;
        RECT 31.460 49.900 31.830 49.910 ;
        RECT 35.305 49.815 36.330 50.075 ;
        RECT 122.065 49.910 123.090 50.170 ;
        RECT 125.940 50.075 126.200 50.425 ;
        RECT 126.565 50.075 126.935 50.085 ;
        RECT 122.065 49.900 122.435 49.910 ;
        RECT 125.910 49.815 126.935 50.075 ;
        RECT 35.960 49.805 36.330 49.815 ;
        RECT 126.565 49.805 126.935 49.815 ;
        RECT 31.460 44.660 31.830 44.670 ;
        RECT 122.065 44.660 122.435 44.670 ;
        RECT 31.460 44.400 32.485 44.660 ;
        RECT 35.960 44.570 36.330 44.580 ;
        RECT 31.460 44.390 31.830 44.400 ;
        RECT 32.195 44.015 32.455 44.400 ;
        RECT 35.305 44.310 36.330 44.570 ;
        RECT 122.065 44.400 123.090 44.660 ;
        RECT 126.565 44.570 126.935 44.580 ;
        RECT 122.065 44.390 122.435 44.400 ;
        RECT 35.335 44.015 35.595 44.310 ;
        RECT 35.960 44.300 36.330 44.310 ;
        RECT 122.800 44.015 123.060 44.400 ;
        RECT 125.910 44.310 126.935 44.570 ;
        RECT 125.940 44.015 126.200 44.310 ;
        RECT 126.565 44.300 126.935 44.310 ;
        RECT 29.785 42.890 127.180 44.015 ;
        RECT 29.785 36.480 30.925 42.890 ;
        RECT 31.460 42.635 31.830 42.645 ;
        RECT 32.195 42.635 32.455 42.890 ;
        RECT 31.460 42.375 32.485 42.635 ;
        RECT 35.335 42.540 35.595 42.890 ;
        RECT 122.065 42.635 122.435 42.645 ;
        RECT 122.800 42.635 123.060 42.890 ;
        RECT 35.960 42.540 36.330 42.550 ;
        RECT 31.460 42.365 31.830 42.375 ;
        RECT 35.305 42.280 36.330 42.540 ;
        RECT 122.065 42.375 123.090 42.635 ;
        RECT 125.940 42.540 126.200 42.890 ;
        RECT 126.565 42.540 126.935 42.550 ;
        RECT 122.065 42.365 122.435 42.375 ;
        RECT 125.910 42.280 126.935 42.540 ;
        RECT 35.960 42.270 36.330 42.280 ;
        RECT 126.565 42.270 126.935 42.280 ;
        RECT 31.460 37.125 31.830 37.135 ;
        RECT 122.065 37.125 122.435 37.135 ;
        RECT 31.460 36.865 32.485 37.125 ;
        RECT 35.960 37.035 36.330 37.045 ;
        RECT 31.460 36.855 31.830 36.865 ;
        RECT 32.195 36.480 32.455 36.865 ;
        RECT 35.305 36.775 36.330 37.035 ;
        RECT 122.065 36.865 123.090 37.125 ;
        RECT 126.565 37.035 126.935 37.045 ;
        RECT 122.065 36.855 122.435 36.865 ;
        RECT 35.335 36.480 35.595 36.775 ;
        RECT 35.960 36.765 36.330 36.775 ;
        RECT 122.800 36.480 123.060 36.865 ;
        RECT 125.910 36.775 126.935 37.035 ;
        RECT 125.940 36.480 126.200 36.775 ;
        RECT 126.565 36.765 126.935 36.775 ;
        RECT 29.785 35.355 127.180 36.480 ;
        RECT 29.785 28.945 30.925 35.355 ;
        RECT 31.460 35.100 31.830 35.110 ;
        RECT 32.195 35.100 32.455 35.355 ;
        RECT 31.460 34.840 32.485 35.100 ;
        RECT 35.335 35.005 35.595 35.355 ;
        RECT 122.065 35.100 122.435 35.110 ;
        RECT 122.800 35.100 123.060 35.355 ;
        RECT 35.960 35.005 36.330 35.015 ;
        RECT 31.460 34.830 31.830 34.840 ;
        RECT 35.305 34.745 36.330 35.005 ;
        RECT 122.065 34.840 123.090 35.100 ;
        RECT 125.940 35.005 126.200 35.355 ;
        RECT 126.565 35.005 126.935 35.015 ;
        RECT 122.065 34.830 122.435 34.840 ;
        RECT 125.910 34.745 126.935 35.005 ;
        RECT 35.960 34.735 36.330 34.745 ;
        RECT 126.565 34.735 126.935 34.745 ;
        RECT 31.460 29.590 31.830 29.600 ;
        RECT 122.065 29.590 122.435 29.600 ;
        RECT 31.460 29.330 32.485 29.590 ;
        RECT 35.960 29.500 36.330 29.510 ;
        RECT 31.460 29.320 31.830 29.330 ;
        RECT 32.195 28.945 32.455 29.330 ;
        RECT 35.305 29.240 36.330 29.500 ;
        RECT 122.065 29.330 123.090 29.590 ;
        RECT 126.565 29.500 126.935 29.510 ;
        RECT 122.065 29.320 122.435 29.330 ;
        RECT 35.335 28.945 35.595 29.240 ;
        RECT 35.960 29.230 36.330 29.240 ;
        RECT 122.800 28.945 123.060 29.330 ;
        RECT 125.910 29.240 126.935 29.500 ;
        RECT 125.940 28.945 126.200 29.240 ;
        RECT 126.565 29.230 126.935 29.240 ;
        RECT 29.785 27.820 127.180 28.945 ;
        RECT 29.785 21.410 30.925 27.820 ;
        RECT 31.460 27.565 31.830 27.575 ;
        RECT 32.195 27.565 32.455 27.820 ;
        RECT 31.460 27.305 32.485 27.565 ;
        RECT 35.335 27.470 35.595 27.820 ;
        RECT 122.065 27.565 122.435 27.575 ;
        RECT 122.800 27.565 123.060 27.820 ;
        RECT 35.960 27.470 36.330 27.480 ;
        RECT 31.460 27.295 31.830 27.305 ;
        RECT 35.305 27.210 36.330 27.470 ;
        RECT 122.065 27.305 123.090 27.565 ;
        RECT 125.940 27.470 126.200 27.820 ;
        RECT 126.565 27.470 126.935 27.480 ;
        RECT 122.065 27.295 122.435 27.305 ;
        RECT 125.910 27.210 126.935 27.470 ;
        RECT 35.960 27.200 36.330 27.210 ;
        RECT 126.565 27.200 126.935 27.210 ;
        RECT 31.460 22.055 31.830 22.065 ;
        RECT 122.065 22.055 122.435 22.065 ;
        RECT 31.460 21.795 32.485 22.055 ;
        RECT 35.960 21.965 36.330 21.975 ;
        RECT 31.460 21.785 31.830 21.795 ;
        RECT 32.195 21.410 32.455 21.795 ;
        RECT 35.305 21.705 36.330 21.965 ;
        RECT 122.065 21.795 123.090 22.055 ;
        RECT 126.565 21.965 126.935 21.975 ;
        RECT 122.065 21.785 122.435 21.795 ;
        RECT 35.335 21.410 35.595 21.705 ;
        RECT 35.960 21.695 36.330 21.705 ;
        RECT 122.800 21.410 123.060 21.795 ;
        RECT 125.910 21.705 126.935 21.965 ;
        RECT 125.940 21.410 126.200 21.705 ;
        RECT 126.565 21.695 126.935 21.705 ;
        RECT 29.785 20.285 127.180 21.410 ;
        RECT 29.785 13.875 30.925 20.285 ;
        RECT 31.460 20.030 31.830 20.040 ;
        RECT 32.195 20.030 32.455 20.285 ;
        RECT 31.460 19.770 32.485 20.030 ;
        RECT 35.335 19.935 35.595 20.285 ;
        RECT 122.065 20.030 122.435 20.040 ;
        RECT 122.800 20.030 123.060 20.285 ;
        RECT 35.960 19.935 36.330 19.945 ;
        RECT 31.460 19.760 31.830 19.770 ;
        RECT 35.305 19.675 36.330 19.935 ;
        RECT 122.065 19.770 123.090 20.030 ;
        RECT 125.940 19.935 126.200 20.285 ;
        RECT 126.565 19.935 126.935 19.945 ;
        RECT 122.065 19.760 122.435 19.770 ;
        RECT 125.910 19.675 126.935 19.935 ;
        RECT 35.960 19.665 36.330 19.675 ;
        RECT 126.565 19.665 126.935 19.675 ;
        RECT 31.460 14.520 31.830 14.530 ;
        RECT 122.065 14.520 122.435 14.530 ;
        RECT 31.460 14.260 32.485 14.520 ;
        RECT 35.960 14.430 36.330 14.440 ;
        RECT 31.460 14.250 31.830 14.260 ;
        RECT 32.195 13.875 32.455 14.260 ;
        RECT 35.305 14.170 36.330 14.430 ;
        RECT 122.065 14.260 123.090 14.520 ;
        RECT 126.565 14.430 126.935 14.440 ;
        RECT 122.065 14.250 122.435 14.260 ;
        RECT 35.335 13.875 35.595 14.170 ;
        RECT 35.960 14.160 36.330 14.170 ;
        RECT 122.800 13.875 123.060 14.260 ;
        RECT 125.910 14.170 126.935 14.430 ;
        RECT 125.940 13.875 126.200 14.170 ;
        RECT 126.565 14.160 126.935 14.170 ;
        RECT 29.785 12.750 127.180 13.875 ;
        RECT 29.785 6.340 30.925 12.750 ;
        RECT 31.460 12.495 31.830 12.505 ;
        RECT 32.195 12.495 32.455 12.750 ;
        RECT 31.460 12.235 32.485 12.495 ;
        RECT 35.335 12.400 35.595 12.750 ;
        RECT 122.065 12.495 122.435 12.505 ;
        RECT 122.800 12.495 123.060 12.750 ;
        RECT 35.960 12.400 36.330 12.410 ;
        RECT 31.460 12.225 31.830 12.235 ;
        RECT 35.305 12.140 36.330 12.400 ;
        RECT 122.065 12.235 123.090 12.495 ;
        RECT 125.940 12.400 126.200 12.750 ;
        RECT 126.565 12.400 126.935 12.410 ;
        RECT 122.065 12.225 122.435 12.235 ;
        RECT 125.910 12.140 126.935 12.400 ;
        RECT 35.960 12.130 36.330 12.140 ;
        RECT 126.565 12.130 126.935 12.140 ;
        RECT 31.460 6.985 31.830 6.995 ;
        RECT 36.785 6.985 37.155 6.995 ;
        RECT 42.120 6.985 42.490 6.995 ;
        RECT 47.445 6.985 47.815 6.995 ;
        RECT 52.780 6.985 53.150 6.995 ;
        RECT 58.105 6.985 58.475 6.995 ;
        RECT 63.440 6.985 63.810 6.995 ;
        RECT 68.765 6.985 69.135 6.995 ;
        RECT 74.100 6.985 74.470 6.995 ;
        RECT 79.425 6.985 79.795 6.995 ;
        RECT 84.760 6.985 85.130 6.995 ;
        RECT 90.085 6.985 90.455 6.995 ;
        RECT 95.420 6.985 95.790 6.995 ;
        RECT 100.745 6.985 101.115 6.995 ;
        RECT 106.080 6.985 106.450 6.995 ;
        RECT 111.405 6.985 111.775 6.995 ;
        RECT 116.740 6.985 117.110 6.995 ;
        RECT 122.065 6.985 122.435 6.995 ;
        RECT 31.460 6.725 32.485 6.985 ;
        RECT 35.960 6.895 36.330 6.905 ;
        RECT 31.460 6.715 31.830 6.725 ;
        RECT 32.195 6.340 32.455 6.725 ;
        RECT 35.305 6.635 36.330 6.895 ;
        RECT 36.785 6.725 37.810 6.985 ;
        RECT 41.285 6.895 41.655 6.905 ;
        RECT 36.785 6.715 37.155 6.725 ;
        RECT 35.335 6.340 35.595 6.635 ;
        RECT 35.960 6.625 36.330 6.635 ;
        RECT 37.520 6.340 37.780 6.725 ;
        RECT 40.630 6.635 41.655 6.895 ;
        RECT 42.120 6.725 43.145 6.985 ;
        RECT 46.620 6.895 46.990 6.905 ;
        RECT 42.120 6.715 42.490 6.725 ;
        RECT 40.660 6.340 40.920 6.635 ;
        RECT 41.285 6.625 41.655 6.635 ;
        RECT 42.855 6.340 43.115 6.725 ;
        RECT 45.965 6.635 46.990 6.895 ;
        RECT 47.445 6.725 48.470 6.985 ;
        RECT 51.945 6.895 52.315 6.905 ;
        RECT 47.445 6.715 47.815 6.725 ;
        RECT 45.995 6.340 46.255 6.635 ;
        RECT 46.620 6.625 46.990 6.635 ;
        RECT 48.180 6.340 48.440 6.725 ;
        RECT 51.290 6.635 52.315 6.895 ;
        RECT 52.780 6.725 53.805 6.985 ;
        RECT 57.280 6.895 57.650 6.905 ;
        RECT 52.780 6.715 53.150 6.725 ;
        RECT 51.320 6.340 51.580 6.635 ;
        RECT 51.945 6.625 52.315 6.635 ;
        RECT 53.515 6.340 53.775 6.725 ;
        RECT 56.625 6.635 57.650 6.895 ;
        RECT 58.105 6.725 59.130 6.985 ;
        RECT 62.605 6.895 62.975 6.905 ;
        RECT 58.105 6.715 58.475 6.725 ;
        RECT 56.655 6.340 56.915 6.635 ;
        RECT 57.280 6.625 57.650 6.635 ;
        RECT 58.840 6.340 59.100 6.725 ;
        RECT 61.950 6.635 62.975 6.895 ;
        RECT 63.440 6.725 64.465 6.985 ;
        RECT 67.940 6.895 68.310 6.905 ;
        RECT 63.440 6.715 63.810 6.725 ;
        RECT 61.980 6.340 62.240 6.635 ;
        RECT 62.605 6.625 62.975 6.635 ;
        RECT 64.175 6.340 64.435 6.725 ;
        RECT 67.285 6.635 68.310 6.895 ;
        RECT 68.765 6.725 69.790 6.985 ;
        RECT 73.265 6.895 73.635 6.905 ;
        RECT 68.765 6.715 69.135 6.725 ;
        RECT 67.315 6.340 67.575 6.635 ;
        RECT 67.940 6.625 68.310 6.635 ;
        RECT 69.500 6.340 69.760 6.725 ;
        RECT 72.610 6.635 73.635 6.895 ;
        RECT 74.100 6.725 75.125 6.985 ;
        RECT 78.600 6.895 78.970 6.905 ;
        RECT 74.100 6.715 74.470 6.725 ;
        RECT 72.640 6.340 72.900 6.635 ;
        RECT 73.265 6.625 73.635 6.635 ;
        RECT 74.835 6.340 75.095 6.725 ;
        RECT 77.945 6.635 78.970 6.895 ;
        RECT 79.425 6.725 80.450 6.985 ;
        RECT 83.925 6.895 84.295 6.905 ;
        RECT 79.425 6.715 79.795 6.725 ;
        RECT 77.975 6.340 78.235 6.635 ;
        RECT 78.600 6.625 78.970 6.635 ;
        RECT 80.160 6.340 80.420 6.725 ;
        RECT 83.270 6.635 84.295 6.895 ;
        RECT 84.760 6.725 85.785 6.985 ;
        RECT 89.260 6.895 89.630 6.905 ;
        RECT 84.760 6.715 85.130 6.725 ;
        RECT 83.300 6.340 83.560 6.635 ;
        RECT 83.925 6.625 84.295 6.635 ;
        RECT 85.495 6.340 85.755 6.725 ;
        RECT 88.605 6.635 89.630 6.895 ;
        RECT 90.085 6.725 91.110 6.985 ;
        RECT 94.585 6.895 94.955 6.905 ;
        RECT 90.085 6.715 90.455 6.725 ;
        RECT 88.635 6.340 88.895 6.635 ;
        RECT 89.260 6.625 89.630 6.635 ;
        RECT 90.820 6.340 91.080 6.725 ;
        RECT 93.930 6.635 94.955 6.895 ;
        RECT 95.420 6.725 96.445 6.985 ;
        RECT 99.920 6.895 100.290 6.905 ;
        RECT 95.420 6.715 95.790 6.725 ;
        RECT 93.960 6.340 94.220 6.635 ;
        RECT 94.585 6.625 94.955 6.635 ;
        RECT 96.155 6.340 96.415 6.725 ;
        RECT 99.265 6.635 100.290 6.895 ;
        RECT 100.745 6.725 101.770 6.985 ;
        RECT 105.245 6.895 105.615 6.905 ;
        RECT 100.745 6.715 101.115 6.725 ;
        RECT 99.295 6.340 99.555 6.635 ;
        RECT 99.920 6.625 100.290 6.635 ;
        RECT 101.480 6.340 101.740 6.725 ;
        RECT 104.590 6.635 105.615 6.895 ;
        RECT 106.080 6.725 107.105 6.985 ;
        RECT 110.580 6.895 110.950 6.905 ;
        RECT 106.080 6.715 106.450 6.725 ;
        RECT 104.620 6.340 104.880 6.635 ;
        RECT 105.245 6.625 105.615 6.635 ;
        RECT 106.815 6.340 107.075 6.725 ;
        RECT 109.925 6.635 110.950 6.895 ;
        RECT 111.405 6.725 112.430 6.985 ;
        RECT 115.905 6.895 116.275 6.905 ;
        RECT 111.405 6.715 111.775 6.725 ;
        RECT 109.955 6.340 110.215 6.635 ;
        RECT 110.580 6.625 110.950 6.635 ;
        RECT 112.140 6.340 112.400 6.725 ;
        RECT 115.250 6.635 116.275 6.895 ;
        RECT 116.740 6.725 117.765 6.985 ;
        RECT 121.240 6.895 121.610 6.905 ;
        RECT 116.740 6.715 117.110 6.725 ;
        RECT 115.280 6.340 115.540 6.635 ;
        RECT 115.905 6.625 116.275 6.635 ;
        RECT 117.475 6.340 117.735 6.725 ;
        RECT 120.585 6.635 121.610 6.895 ;
        RECT 122.065 6.725 123.090 6.985 ;
        RECT 126.565 6.895 126.935 6.905 ;
        RECT 122.065 6.715 122.435 6.725 ;
        RECT 120.615 6.340 120.875 6.635 ;
        RECT 121.240 6.625 121.610 6.635 ;
        RECT 122.800 6.340 123.060 6.725 ;
        RECT 125.910 6.635 126.935 6.895 ;
        RECT 125.940 6.340 126.200 6.635 ;
        RECT 126.565 6.625 126.935 6.635 ;
        RECT 29.785 5.215 127.180 6.340 ;
        RECT 29.785 1.085 30.925 5.215 ;
        RECT 31.460 4.960 31.830 4.970 ;
        RECT 32.195 4.960 32.455 5.215 ;
        RECT 31.460 4.700 32.485 4.960 ;
        RECT 35.335 4.865 35.595 5.215 ;
        RECT 36.785 4.960 37.155 4.970 ;
        RECT 37.520 4.960 37.780 5.215 ;
        RECT 35.960 4.865 36.330 4.875 ;
        RECT 31.460 4.690 31.830 4.700 ;
        RECT 35.305 4.605 36.330 4.865 ;
        RECT 36.785 4.700 37.810 4.960 ;
        RECT 40.660 4.865 40.920 5.215 ;
        RECT 42.120 4.960 42.490 4.970 ;
        RECT 42.855 4.960 43.115 5.215 ;
        RECT 41.285 4.865 41.655 4.875 ;
        RECT 36.785 4.690 37.155 4.700 ;
        RECT 40.630 4.605 41.655 4.865 ;
        RECT 42.120 4.700 43.145 4.960 ;
        RECT 45.995 4.865 46.255 5.215 ;
        RECT 47.445 4.960 47.815 4.970 ;
        RECT 48.180 4.960 48.440 5.215 ;
        RECT 46.620 4.865 46.990 4.875 ;
        RECT 42.120 4.690 42.490 4.700 ;
        RECT 45.965 4.605 46.990 4.865 ;
        RECT 47.445 4.700 48.470 4.960 ;
        RECT 51.320 4.865 51.580 5.215 ;
        RECT 52.780 4.960 53.150 4.970 ;
        RECT 53.515 4.960 53.775 5.215 ;
        RECT 51.945 4.865 52.315 4.875 ;
        RECT 47.445 4.690 47.815 4.700 ;
        RECT 51.290 4.605 52.315 4.865 ;
        RECT 52.780 4.700 53.805 4.960 ;
        RECT 56.655 4.865 56.915 5.215 ;
        RECT 58.105 4.960 58.475 4.970 ;
        RECT 58.840 4.960 59.100 5.215 ;
        RECT 57.280 4.865 57.650 4.875 ;
        RECT 52.780 4.690 53.150 4.700 ;
        RECT 56.625 4.605 57.650 4.865 ;
        RECT 58.105 4.700 59.130 4.960 ;
        RECT 61.980 4.865 62.240 5.215 ;
        RECT 63.440 4.960 63.810 4.970 ;
        RECT 64.175 4.960 64.435 5.215 ;
        RECT 62.605 4.865 62.975 4.875 ;
        RECT 58.105 4.690 58.475 4.700 ;
        RECT 61.950 4.605 62.975 4.865 ;
        RECT 63.440 4.700 64.465 4.960 ;
        RECT 67.315 4.865 67.575 5.215 ;
        RECT 68.765 4.960 69.135 4.970 ;
        RECT 69.500 4.960 69.760 5.215 ;
        RECT 67.940 4.865 68.310 4.875 ;
        RECT 63.440 4.690 63.810 4.700 ;
        RECT 67.285 4.605 68.310 4.865 ;
        RECT 68.765 4.700 69.790 4.960 ;
        RECT 72.640 4.865 72.900 5.215 ;
        RECT 74.100 4.960 74.470 4.970 ;
        RECT 74.835 4.960 75.095 5.215 ;
        RECT 73.265 4.865 73.635 4.875 ;
        RECT 68.765 4.690 69.135 4.700 ;
        RECT 72.610 4.605 73.635 4.865 ;
        RECT 74.100 4.700 75.125 4.960 ;
        RECT 77.975 4.865 78.235 5.215 ;
        RECT 79.425 4.960 79.795 4.970 ;
        RECT 80.160 4.960 80.420 5.215 ;
        RECT 78.600 4.865 78.970 4.875 ;
        RECT 74.100 4.690 74.470 4.700 ;
        RECT 77.945 4.605 78.970 4.865 ;
        RECT 79.425 4.700 80.450 4.960 ;
        RECT 83.300 4.865 83.560 5.215 ;
        RECT 84.760 4.960 85.130 4.970 ;
        RECT 85.495 4.960 85.755 5.215 ;
        RECT 83.925 4.865 84.295 4.875 ;
        RECT 79.425 4.690 79.795 4.700 ;
        RECT 83.270 4.605 84.295 4.865 ;
        RECT 84.760 4.700 85.785 4.960 ;
        RECT 88.635 4.865 88.895 5.215 ;
        RECT 90.085 4.960 90.455 4.970 ;
        RECT 90.820 4.960 91.080 5.215 ;
        RECT 89.260 4.865 89.630 4.875 ;
        RECT 84.760 4.690 85.130 4.700 ;
        RECT 88.605 4.605 89.630 4.865 ;
        RECT 90.085 4.700 91.110 4.960 ;
        RECT 93.960 4.865 94.220 5.215 ;
        RECT 95.420 4.960 95.790 4.970 ;
        RECT 96.155 4.960 96.415 5.215 ;
        RECT 94.585 4.865 94.955 4.875 ;
        RECT 90.085 4.690 90.455 4.700 ;
        RECT 93.930 4.605 94.955 4.865 ;
        RECT 95.420 4.700 96.445 4.960 ;
        RECT 99.295 4.865 99.555 5.215 ;
        RECT 100.745 4.960 101.115 4.970 ;
        RECT 101.480 4.960 101.740 5.215 ;
        RECT 99.920 4.865 100.290 4.875 ;
        RECT 95.420 4.690 95.790 4.700 ;
        RECT 99.265 4.605 100.290 4.865 ;
        RECT 100.745 4.700 101.770 4.960 ;
        RECT 104.620 4.865 104.880 5.215 ;
        RECT 106.080 4.960 106.450 4.970 ;
        RECT 106.815 4.960 107.075 5.215 ;
        RECT 105.245 4.865 105.615 4.875 ;
        RECT 100.745 4.690 101.115 4.700 ;
        RECT 104.590 4.605 105.615 4.865 ;
        RECT 106.080 4.700 107.105 4.960 ;
        RECT 109.955 4.865 110.215 5.215 ;
        RECT 111.405 4.960 111.775 4.970 ;
        RECT 112.140 4.960 112.400 5.215 ;
        RECT 110.580 4.865 110.950 4.875 ;
        RECT 106.080 4.690 106.450 4.700 ;
        RECT 109.925 4.605 110.950 4.865 ;
        RECT 111.405 4.700 112.430 4.960 ;
        RECT 115.280 4.865 115.540 5.215 ;
        RECT 116.740 4.960 117.110 4.970 ;
        RECT 117.475 4.960 117.735 5.215 ;
        RECT 115.905 4.865 116.275 4.875 ;
        RECT 111.405 4.690 111.775 4.700 ;
        RECT 115.250 4.605 116.275 4.865 ;
        RECT 116.740 4.700 117.765 4.960 ;
        RECT 120.615 4.865 120.875 5.215 ;
        RECT 122.065 4.960 122.435 4.970 ;
        RECT 122.800 4.960 123.060 5.215 ;
        RECT 121.240 4.865 121.610 4.875 ;
        RECT 116.740 4.690 117.110 4.700 ;
        RECT 120.585 4.605 121.610 4.865 ;
        RECT 122.065 4.700 123.090 4.960 ;
        RECT 125.940 4.865 126.200 5.215 ;
        RECT 126.565 4.865 126.935 4.875 ;
        RECT 122.065 4.690 122.435 4.700 ;
        RECT 125.910 4.605 126.935 4.865 ;
        RECT 35.960 4.595 36.330 4.605 ;
        RECT 41.285 4.595 41.655 4.605 ;
        RECT 46.620 4.595 46.990 4.605 ;
        RECT 51.945 4.595 52.315 4.605 ;
        RECT 57.280 4.595 57.650 4.605 ;
        RECT 62.605 4.595 62.975 4.605 ;
        RECT 67.940 4.595 68.310 4.605 ;
        RECT 73.265 4.595 73.635 4.605 ;
        RECT 78.600 4.595 78.970 4.605 ;
        RECT 83.925 4.595 84.295 4.605 ;
        RECT 89.260 4.595 89.630 4.605 ;
        RECT 94.585 4.595 94.955 4.605 ;
        RECT 99.920 4.595 100.290 4.605 ;
        RECT 105.245 4.595 105.615 4.605 ;
        RECT 110.580 4.595 110.950 4.605 ;
        RECT 115.905 4.595 116.275 4.605 ;
        RECT 121.240 4.595 121.610 4.605 ;
        RECT 126.565 4.595 126.935 4.605 ;
      LAYER met3 ;
        RECT 26.760 83.390 74.685 84.455 ;
        RECT 26.760 83.090 75.720 83.390 ;
        RECT 26.760 81.830 74.685 83.090 ;
        RECT 26.760 79.635 30.970 81.830 ;
        RECT -1.000 76.265 30.970 79.635 ;
        RECT 29.740 70.565 30.970 76.265 ;
        RECT 31.480 74.420 31.810 75.175 ;
        RECT 35.980 74.020 36.310 74.770 ;
        RECT 36.805 74.420 37.135 75.175 ;
        RECT 41.305 74.020 41.635 74.770 ;
        RECT 42.140 74.420 42.470 75.175 ;
        RECT 46.640 74.020 46.970 74.770 ;
        RECT 47.465 74.420 47.795 75.175 ;
        RECT 51.965 74.020 52.295 74.770 ;
        RECT 52.800 74.420 53.130 75.175 ;
        RECT 57.300 74.020 57.630 74.770 ;
        RECT 58.125 74.420 58.455 75.175 ;
        RECT 62.625 74.020 62.955 74.770 ;
        RECT 63.460 74.420 63.790 75.175 ;
        RECT 67.960 74.020 68.290 74.770 ;
        RECT 68.785 74.420 69.115 75.175 ;
        RECT 73.285 74.020 73.615 74.770 ;
        RECT 74.120 74.420 74.450 75.175 ;
        RECT 31.480 72.455 31.810 73.205 ;
        RECT 35.980 71.970 36.310 72.730 ;
        RECT 36.805 72.455 37.135 73.205 ;
        RECT 41.305 71.970 41.635 72.730 ;
        RECT 42.140 72.455 42.470 73.205 ;
        RECT 46.640 71.970 46.970 72.730 ;
        RECT 47.465 72.455 47.795 73.205 ;
        RECT 51.965 71.970 52.295 72.730 ;
        RECT 52.800 72.455 53.130 73.205 ;
        RECT 57.300 71.970 57.630 72.730 ;
        RECT 58.125 72.455 58.455 73.205 ;
        RECT 62.625 71.970 62.955 72.730 ;
        RECT 63.460 72.455 63.790 73.205 ;
        RECT 67.960 71.970 68.290 72.730 ;
        RECT 68.785 72.455 69.115 73.205 ;
        RECT 73.285 71.970 73.615 72.730 ;
        RECT 74.120 72.455 74.450 73.205 ;
        RECT 75.420 68.495 75.720 83.090 ;
        RECT 118.060 78.530 118.770 80.280 ;
        RECT 78.620 74.020 78.950 74.770 ;
        RECT 79.445 74.420 79.775 75.175 ;
        RECT 83.945 74.020 84.275 74.770 ;
        RECT 84.780 74.420 85.110 75.175 ;
        RECT 89.280 74.020 89.610 74.770 ;
        RECT 90.105 74.420 90.435 75.175 ;
        RECT 94.605 74.020 94.935 74.770 ;
        RECT 95.440 74.420 95.770 75.175 ;
        RECT 99.940 74.020 100.270 74.770 ;
        RECT 100.765 74.420 101.095 75.175 ;
        RECT 105.265 74.020 105.595 74.770 ;
        RECT 106.100 74.420 106.430 75.175 ;
        RECT 110.600 74.020 110.930 74.770 ;
        RECT 111.425 74.420 111.755 75.175 ;
        RECT 115.925 74.020 116.255 74.770 ;
        RECT 116.760 74.420 117.090 75.175 ;
        RECT 78.620 71.970 78.950 72.730 ;
        RECT 79.445 72.455 79.775 73.205 ;
        RECT 83.945 71.970 84.275 72.730 ;
        RECT 84.780 72.455 85.110 73.205 ;
        RECT 89.280 71.970 89.610 72.730 ;
        RECT 90.105 72.455 90.435 73.205 ;
        RECT 94.605 71.970 94.935 72.730 ;
        RECT 95.440 72.455 95.770 73.205 ;
        RECT 99.940 71.970 100.270 72.730 ;
        RECT 100.765 72.455 101.095 73.205 ;
        RECT 105.265 71.970 105.595 72.730 ;
        RECT 106.100 72.455 106.430 73.205 ;
        RECT 110.600 71.970 110.930 72.730 ;
        RECT 111.425 72.455 111.755 73.205 ;
        RECT 115.925 71.970 116.255 72.730 ;
        RECT 116.760 72.455 117.090 73.205 ;
        RECT 118.060 68.495 118.360 78.530 ;
        RECT 121.260 74.020 121.590 74.770 ;
        RECT 122.085 74.420 122.415 75.175 ;
        RECT 126.585 74.020 126.915 74.770 ;
        RECT 121.260 71.970 121.590 72.730 ;
        RECT 122.085 72.455 122.415 73.205 ;
        RECT 126.585 71.970 126.915 72.730 ;
        RECT 74.120 68.195 75.720 68.495 ;
        RECT 116.760 68.195 118.360 68.495 ;
        RECT 31.480 66.885 31.810 67.640 ;
        RECT 35.980 66.485 36.310 67.235 ;
        RECT 74.120 66.935 74.450 68.195 ;
        RECT 116.760 66.935 117.090 68.195 ;
        RECT 122.085 66.885 122.415 67.640 ;
        RECT 126.585 66.485 126.915 67.235 ;
        RECT 31.480 64.920 31.810 65.670 ;
        RECT 35.980 64.435 36.310 65.195 ;
        RECT 122.085 64.920 122.415 65.670 ;
        RECT 126.585 64.435 126.915 65.195 ;
        RECT 31.480 59.350 31.810 60.105 ;
        RECT 35.980 58.950 36.310 59.700 ;
        RECT 122.085 59.350 122.415 60.105 ;
        RECT 126.585 58.950 126.915 59.700 ;
        RECT 31.480 57.385 31.810 58.135 ;
        RECT 35.980 56.900 36.310 57.660 ;
        RECT 122.085 57.385 122.415 58.135 ;
        RECT 126.585 56.900 126.915 57.660 ;
        RECT 31.480 51.815 31.810 52.570 ;
        RECT 35.980 51.415 36.310 52.165 ;
        RECT 122.085 51.815 122.415 52.570 ;
        RECT 126.585 51.415 126.915 52.165 ;
        RECT 31.480 49.850 31.810 50.600 ;
        RECT 35.980 49.365 36.310 50.125 ;
        RECT 122.085 49.850 122.415 50.600 ;
        RECT 126.585 49.365 126.915 50.125 ;
        RECT 31.480 44.280 31.810 45.035 ;
        RECT 35.980 43.880 36.310 44.630 ;
        RECT 122.085 44.280 122.415 45.035 ;
        RECT 126.585 43.880 126.915 44.630 ;
        RECT 31.480 42.315 31.810 43.065 ;
        RECT 35.980 41.830 36.310 42.590 ;
        RECT 122.085 42.315 122.415 43.065 ;
        RECT 126.585 41.830 126.915 42.590 ;
        RECT 31.480 36.745 31.810 37.500 ;
        RECT 35.980 36.345 36.310 37.095 ;
        RECT 122.085 36.745 122.415 37.500 ;
        RECT 126.585 36.345 126.915 37.095 ;
        RECT 31.480 34.780 31.810 35.530 ;
        RECT 35.980 34.295 36.310 35.055 ;
        RECT 122.085 34.780 122.415 35.530 ;
        RECT 126.585 34.295 126.915 35.055 ;
        RECT 31.480 29.210 31.810 29.965 ;
        RECT 35.980 28.810 36.310 29.560 ;
        RECT 122.085 29.210 122.415 29.965 ;
        RECT 126.585 28.810 126.915 29.560 ;
        RECT 31.480 27.245 31.810 27.995 ;
        RECT 35.980 26.760 36.310 27.520 ;
        RECT 122.085 27.245 122.415 27.995 ;
        RECT 126.585 26.760 126.915 27.520 ;
        RECT 31.480 21.675 31.810 22.430 ;
        RECT 35.980 21.275 36.310 22.025 ;
        RECT 122.085 21.675 122.415 22.430 ;
        RECT 126.585 21.275 126.915 22.025 ;
        RECT 31.480 19.710 31.810 20.460 ;
        RECT 35.980 19.225 36.310 19.985 ;
        RECT 122.085 19.710 122.415 20.460 ;
        RECT 126.585 19.225 126.915 19.985 ;
        RECT 31.480 14.140 31.810 14.895 ;
        RECT 35.980 13.740 36.310 14.490 ;
        RECT 122.085 14.140 122.415 14.895 ;
        RECT 126.585 13.740 126.915 14.490 ;
        RECT 31.480 12.175 31.810 12.925 ;
        RECT 35.980 11.690 36.310 12.450 ;
        RECT 122.085 12.175 122.415 12.925 ;
        RECT 126.585 11.690 126.915 12.450 ;
        RECT 31.480 6.605 31.810 7.360 ;
        RECT 35.980 6.205 36.310 6.955 ;
        RECT 36.805 6.605 37.135 7.360 ;
        RECT 41.305 6.205 41.635 6.955 ;
        RECT 42.140 6.605 42.470 7.360 ;
        RECT 46.640 6.205 46.970 6.955 ;
        RECT 47.465 6.605 47.795 7.360 ;
        RECT 51.965 6.205 52.295 6.955 ;
        RECT 52.800 6.605 53.130 7.360 ;
        RECT 57.300 6.205 57.630 6.955 ;
        RECT 58.125 6.605 58.455 7.360 ;
        RECT 62.625 6.205 62.955 6.955 ;
        RECT 63.460 6.605 63.790 7.360 ;
        RECT 67.960 6.205 68.290 6.955 ;
        RECT 68.785 6.605 69.115 7.360 ;
        RECT 73.285 6.205 73.615 6.955 ;
        RECT 74.120 6.605 74.450 7.360 ;
        RECT 78.620 6.205 78.950 6.955 ;
        RECT 79.445 6.605 79.775 7.360 ;
        RECT 83.945 6.205 84.275 6.955 ;
        RECT 84.780 6.605 85.110 7.360 ;
        RECT 89.280 6.205 89.610 6.955 ;
        RECT 90.105 6.605 90.435 7.360 ;
        RECT 94.605 6.205 94.935 6.955 ;
        RECT 95.440 6.605 95.770 7.360 ;
        RECT 99.940 6.205 100.270 6.955 ;
        RECT 100.765 6.605 101.095 7.360 ;
        RECT 105.265 6.205 105.595 6.955 ;
        RECT 106.100 6.605 106.430 7.360 ;
        RECT 110.600 6.205 110.930 6.955 ;
        RECT 111.425 6.605 111.755 7.360 ;
        RECT 115.925 6.205 116.255 6.955 ;
        RECT 116.760 6.605 117.090 7.360 ;
        RECT 121.260 6.205 121.590 6.955 ;
        RECT 122.085 6.605 122.415 7.360 ;
        RECT 31.480 4.640 31.810 5.390 ;
        RECT 35.980 4.155 36.310 4.915 ;
        RECT 36.805 4.640 37.135 5.390 ;
        RECT 41.305 4.155 41.635 4.915 ;
        RECT 42.140 4.640 42.470 5.390 ;
        RECT 46.640 4.155 46.970 4.915 ;
        RECT 47.465 4.640 47.795 5.390 ;
        RECT 51.965 4.155 52.295 4.915 ;
        RECT 52.800 4.640 53.130 5.390 ;
        RECT 57.300 4.155 57.630 4.915 ;
        RECT 58.125 4.640 58.455 5.390 ;
        RECT 62.625 4.155 62.955 4.915 ;
        RECT 63.460 4.640 63.790 5.390 ;
        RECT 67.960 4.155 68.290 4.915 ;
        RECT 68.785 4.640 69.115 5.390 ;
        RECT 73.285 4.155 73.615 4.915 ;
        RECT 74.120 4.640 74.450 5.390 ;
        RECT 78.620 4.155 78.950 4.915 ;
        RECT 79.445 4.640 79.775 5.390 ;
        RECT 83.945 4.155 84.275 4.915 ;
        RECT 84.780 4.640 85.110 5.390 ;
        RECT 89.280 4.155 89.610 4.915 ;
        RECT 90.105 4.640 90.435 5.390 ;
        RECT 94.605 4.155 94.935 4.915 ;
        RECT 95.440 4.640 95.770 5.390 ;
        RECT 99.940 4.155 100.270 4.915 ;
        RECT 100.765 4.640 101.095 5.390 ;
        RECT 105.265 4.155 105.595 4.915 ;
        RECT 106.100 4.640 106.430 5.390 ;
        RECT 110.600 4.155 110.930 4.915 ;
        RECT 111.425 4.640 111.755 5.390 ;
        RECT 115.925 4.155 116.255 4.915 ;
        RECT 116.760 4.640 117.090 5.390 ;
        RECT 121.260 4.155 121.590 4.915 ;
        RECT 122.085 4.640 122.415 5.390 ;
        RECT 124.185 2.280 125.195 6.340 ;
        RECT 126.585 6.205 126.915 6.955 ;
        RECT 126.585 4.155 126.915 4.915 ;
        RECT 124.185 0.330 129.370 2.280 ;
        RECT 124.185 -0.020 125.985 0.330 ;
      LAYER met4 ;
        RECT 26.755 78.415 129.375 80.545 ;
        RECT 31.480 75.070 31.810 75.085 ;
        RECT 36.805 75.070 37.135 75.085 ;
        RECT 42.140 75.070 42.470 75.085 ;
        RECT 47.465 75.070 47.795 75.085 ;
        RECT 52.800 75.070 53.130 75.085 ;
        RECT 58.125 75.070 58.455 75.085 ;
        RECT 63.460 75.070 63.790 75.085 ;
        RECT 68.785 75.070 69.115 75.085 ;
        RECT 74.120 75.070 74.450 75.085 ;
        RECT 79.445 75.070 79.775 75.085 ;
        RECT 84.780 75.070 85.110 75.085 ;
        RECT 90.105 75.070 90.435 75.085 ;
        RECT 95.440 75.070 95.770 75.085 ;
        RECT 100.765 75.070 101.095 75.085 ;
        RECT 106.100 75.070 106.430 75.085 ;
        RECT 111.425 75.070 111.755 75.085 ;
        RECT 116.760 75.070 117.090 75.085 ;
        RECT 122.085 75.070 122.415 75.085 ;
        RECT 31.240 74.770 127.180 75.070 ;
        RECT 31.480 74.755 31.810 74.770 ;
        RECT 36.805 74.755 37.135 74.770 ;
        RECT 42.140 74.755 42.470 74.770 ;
        RECT 47.465 74.755 47.795 74.770 ;
        RECT 52.800 74.755 53.130 74.770 ;
        RECT 58.125 74.755 58.455 74.770 ;
        RECT 63.460 74.755 63.790 74.770 ;
        RECT 68.785 74.755 69.115 74.770 ;
        RECT 74.120 74.755 74.450 74.770 ;
        RECT 79.445 74.755 79.775 74.770 ;
        RECT 84.780 74.755 85.110 74.770 ;
        RECT 90.105 74.755 90.435 74.770 ;
        RECT 95.440 74.755 95.770 74.770 ;
        RECT 100.765 74.755 101.095 74.770 ;
        RECT 106.100 74.755 106.430 74.770 ;
        RECT 111.425 74.755 111.755 74.770 ;
        RECT 116.760 74.755 117.090 74.770 ;
        RECT 122.085 74.755 122.415 74.770 ;
        RECT 35.980 74.425 36.310 74.440 ;
        RECT 41.305 74.425 41.635 74.440 ;
        RECT 46.640 74.425 46.970 74.440 ;
        RECT 51.965 74.425 52.295 74.440 ;
        RECT 57.300 74.425 57.630 74.440 ;
        RECT 62.625 74.425 62.955 74.440 ;
        RECT 67.960 74.425 68.290 74.440 ;
        RECT 73.285 74.425 73.615 74.440 ;
        RECT 78.620 74.425 78.950 74.440 ;
        RECT 83.945 74.425 84.275 74.440 ;
        RECT 89.280 74.425 89.610 74.440 ;
        RECT 94.605 74.425 94.935 74.440 ;
        RECT 99.940 74.425 100.270 74.440 ;
        RECT 105.265 74.425 105.595 74.440 ;
        RECT 110.600 74.425 110.930 74.440 ;
        RECT 115.925 74.425 116.255 74.440 ;
        RECT 121.260 74.425 121.590 74.440 ;
        RECT 126.585 74.425 126.915 74.440 ;
        RECT 31.240 74.125 127.180 74.425 ;
        RECT 35.980 74.110 36.310 74.125 ;
        RECT 41.305 74.110 41.635 74.125 ;
        RECT 46.640 74.110 46.970 74.125 ;
        RECT 51.965 74.110 52.295 74.125 ;
        RECT 57.300 74.110 57.630 74.125 ;
        RECT 62.625 74.110 62.955 74.125 ;
        RECT 67.960 74.110 68.290 74.125 ;
        RECT 73.285 74.110 73.615 74.125 ;
        RECT 78.620 74.110 78.950 74.125 ;
        RECT 83.945 74.110 84.275 74.125 ;
        RECT 89.280 74.110 89.610 74.125 ;
        RECT 94.605 74.110 94.935 74.125 ;
        RECT 99.940 74.110 100.270 74.125 ;
        RECT 105.265 74.110 105.595 74.125 ;
        RECT 110.600 74.110 110.930 74.125 ;
        RECT 115.925 74.110 116.255 74.125 ;
        RECT 121.260 74.110 121.590 74.125 ;
        RECT 126.585 74.110 126.915 74.125 ;
        RECT 31.480 73.090 31.810 73.105 ;
        RECT 36.805 73.090 37.135 73.105 ;
        RECT 42.140 73.090 42.470 73.105 ;
        RECT 47.465 73.090 47.795 73.105 ;
        RECT 52.800 73.090 53.130 73.105 ;
        RECT 58.125 73.090 58.455 73.105 ;
        RECT 63.460 73.090 63.790 73.105 ;
        RECT 68.785 73.090 69.115 73.105 ;
        RECT 74.120 73.090 74.450 73.105 ;
        RECT 79.445 73.090 79.775 73.105 ;
        RECT 84.780 73.090 85.110 73.105 ;
        RECT 90.105 73.090 90.435 73.105 ;
        RECT 95.440 73.090 95.770 73.105 ;
        RECT 100.765 73.090 101.095 73.105 ;
        RECT 106.100 73.090 106.430 73.105 ;
        RECT 111.425 73.090 111.755 73.105 ;
        RECT 116.760 73.090 117.090 73.105 ;
        RECT 122.085 73.090 122.415 73.105 ;
        RECT 31.240 72.790 127.180 73.090 ;
        RECT 31.480 72.775 31.810 72.790 ;
        RECT 36.805 72.775 37.135 72.790 ;
        RECT 42.140 72.775 42.470 72.790 ;
        RECT 47.465 72.775 47.795 72.790 ;
        RECT 52.800 72.775 53.130 72.790 ;
        RECT 58.125 72.775 58.455 72.790 ;
        RECT 63.460 72.775 63.790 72.790 ;
        RECT 68.785 72.775 69.115 72.790 ;
        RECT 74.120 72.775 74.450 72.790 ;
        RECT 79.445 72.775 79.775 72.790 ;
        RECT 84.780 72.775 85.110 72.790 ;
        RECT 90.105 72.775 90.435 72.790 ;
        RECT 95.440 72.775 95.770 72.790 ;
        RECT 100.765 72.775 101.095 72.790 ;
        RECT 106.100 72.775 106.430 72.790 ;
        RECT 111.425 72.775 111.755 72.790 ;
        RECT 116.760 72.775 117.090 72.790 ;
        RECT 122.085 72.775 122.415 72.790 ;
        RECT 35.980 72.445 36.310 72.460 ;
        RECT 41.305 72.445 41.635 72.460 ;
        RECT 46.640 72.445 46.970 72.460 ;
        RECT 51.965 72.445 52.295 72.460 ;
        RECT 57.300 72.445 57.630 72.460 ;
        RECT 62.625 72.445 62.955 72.460 ;
        RECT 67.960 72.445 68.290 72.460 ;
        RECT 73.285 72.445 73.615 72.460 ;
        RECT 78.620 72.445 78.950 72.460 ;
        RECT 83.945 72.445 84.275 72.460 ;
        RECT 89.280 72.445 89.610 72.460 ;
        RECT 94.605 72.445 94.935 72.460 ;
        RECT 99.940 72.445 100.270 72.460 ;
        RECT 105.265 72.445 105.595 72.460 ;
        RECT 110.600 72.445 110.930 72.460 ;
        RECT 115.925 72.445 116.255 72.460 ;
        RECT 121.260 72.445 121.590 72.460 ;
        RECT 126.585 72.445 126.915 72.460 ;
        RECT 31.240 72.145 127.180 72.445 ;
        RECT 35.980 72.130 36.310 72.145 ;
        RECT 41.305 72.130 41.635 72.145 ;
        RECT 46.640 72.130 46.970 72.145 ;
        RECT 51.965 72.130 52.295 72.145 ;
        RECT 57.300 72.130 57.630 72.145 ;
        RECT 62.625 72.130 62.955 72.145 ;
        RECT 67.960 72.130 68.290 72.145 ;
        RECT 73.285 72.130 73.615 72.145 ;
        RECT 78.620 72.130 78.950 72.145 ;
        RECT 83.945 72.130 84.275 72.145 ;
        RECT 89.280 72.130 89.610 72.145 ;
        RECT 94.605 72.130 94.935 72.145 ;
        RECT 99.940 72.130 100.270 72.145 ;
        RECT 105.265 72.130 105.595 72.145 ;
        RECT 110.600 72.130 110.930 72.145 ;
        RECT 115.925 72.130 116.255 72.145 ;
        RECT 121.260 72.130 121.590 72.145 ;
        RECT 126.585 72.130 126.915 72.145 ;
        RECT 31.480 7.255 31.810 7.270 ;
        RECT 36.805 7.255 37.135 7.270 ;
        RECT 42.140 7.255 42.470 7.270 ;
        RECT 47.465 7.255 47.795 7.270 ;
        RECT 52.800 7.255 53.130 7.270 ;
        RECT 58.125 7.255 58.455 7.270 ;
        RECT 63.460 7.255 63.790 7.270 ;
        RECT 68.785 7.255 69.115 7.270 ;
        RECT 74.120 7.255 74.450 7.270 ;
        RECT 79.445 7.255 79.775 7.270 ;
        RECT 84.780 7.255 85.110 7.270 ;
        RECT 90.105 7.255 90.435 7.270 ;
        RECT 95.440 7.255 95.770 7.270 ;
        RECT 100.765 7.255 101.095 7.270 ;
        RECT 106.100 7.255 106.430 7.270 ;
        RECT 111.425 7.255 111.755 7.270 ;
        RECT 116.760 7.255 117.090 7.270 ;
        RECT 122.085 7.255 122.415 7.270 ;
        RECT 31.240 6.955 127.180 7.255 ;
        RECT 31.480 6.940 31.810 6.955 ;
        RECT 36.805 6.940 37.135 6.955 ;
        RECT 42.140 6.940 42.470 6.955 ;
        RECT 47.465 6.940 47.795 6.955 ;
        RECT 52.800 6.940 53.130 6.955 ;
        RECT 58.125 6.940 58.455 6.955 ;
        RECT 63.460 6.940 63.790 6.955 ;
        RECT 68.785 6.940 69.115 6.955 ;
        RECT 74.120 6.940 74.450 6.955 ;
        RECT 79.445 6.940 79.775 6.955 ;
        RECT 84.780 6.940 85.110 6.955 ;
        RECT 90.105 6.940 90.435 6.955 ;
        RECT 95.440 6.940 95.770 6.955 ;
        RECT 100.765 6.940 101.095 6.955 ;
        RECT 106.100 6.940 106.430 6.955 ;
        RECT 111.425 6.940 111.755 6.955 ;
        RECT 116.760 6.940 117.090 6.955 ;
        RECT 122.085 6.940 122.415 6.955 ;
        RECT 35.980 6.610 36.310 6.625 ;
        RECT 41.305 6.610 41.635 6.625 ;
        RECT 46.640 6.610 46.970 6.625 ;
        RECT 51.965 6.610 52.295 6.625 ;
        RECT 57.300 6.610 57.630 6.625 ;
        RECT 62.625 6.610 62.955 6.625 ;
        RECT 67.960 6.610 68.290 6.625 ;
        RECT 73.285 6.610 73.615 6.625 ;
        RECT 78.620 6.610 78.950 6.625 ;
        RECT 83.945 6.610 84.275 6.625 ;
        RECT 89.280 6.610 89.610 6.625 ;
        RECT 94.605 6.610 94.935 6.625 ;
        RECT 99.940 6.610 100.270 6.625 ;
        RECT 105.265 6.610 105.595 6.625 ;
        RECT 110.600 6.610 110.930 6.625 ;
        RECT 115.925 6.610 116.255 6.625 ;
        RECT 121.260 6.610 121.590 6.625 ;
        RECT 126.585 6.610 126.915 6.625 ;
        RECT 31.240 6.310 127.180 6.610 ;
        RECT 35.980 6.295 36.310 6.310 ;
        RECT 41.305 6.295 41.635 6.310 ;
        RECT 46.640 6.295 46.970 6.310 ;
        RECT 51.965 6.295 52.295 6.310 ;
        RECT 57.300 6.295 57.630 6.310 ;
        RECT 62.625 6.295 62.955 6.310 ;
        RECT 67.960 6.295 68.290 6.310 ;
        RECT 73.285 6.295 73.615 6.310 ;
        RECT 78.620 6.295 78.950 6.310 ;
        RECT 83.945 6.295 84.275 6.310 ;
        RECT 89.280 6.295 89.610 6.310 ;
        RECT 94.605 6.295 94.935 6.310 ;
        RECT 99.940 6.295 100.270 6.310 ;
        RECT 105.265 6.295 105.595 6.310 ;
        RECT 110.600 6.295 110.930 6.310 ;
        RECT 115.925 6.295 116.255 6.310 ;
        RECT 121.260 6.295 121.590 6.310 ;
        RECT 126.585 6.295 126.915 6.310 ;
        RECT 31.480 5.275 31.810 5.290 ;
        RECT 36.805 5.275 37.135 5.290 ;
        RECT 42.140 5.275 42.470 5.290 ;
        RECT 47.465 5.275 47.795 5.290 ;
        RECT 52.800 5.275 53.130 5.290 ;
        RECT 58.125 5.275 58.455 5.290 ;
        RECT 63.460 5.275 63.790 5.290 ;
        RECT 68.785 5.275 69.115 5.290 ;
        RECT 74.120 5.275 74.450 5.290 ;
        RECT 79.445 5.275 79.775 5.290 ;
        RECT 84.780 5.275 85.110 5.290 ;
        RECT 90.105 5.275 90.435 5.290 ;
        RECT 95.440 5.275 95.770 5.290 ;
        RECT 100.765 5.275 101.095 5.290 ;
        RECT 106.100 5.275 106.430 5.290 ;
        RECT 111.425 5.275 111.755 5.290 ;
        RECT 116.760 5.275 117.090 5.290 ;
        RECT 122.085 5.275 122.415 5.290 ;
        RECT 31.240 4.975 127.180 5.275 ;
        RECT 31.480 4.960 31.810 4.975 ;
        RECT 36.805 4.960 37.135 4.975 ;
        RECT 42.140 4.960 42.470 4.975 ;
        RECT 47.465 4.960 47.795 4.975 ;
        RECT 52.800 4.960 53.130 4.975 ;
        RECT 58.125 4.960 58.455 4.975 ;
        RECT 63.460 4.960 63.790 4.975 ;
        RECT 68.785 4.960 69.115 4.975 ;
        RECT 74.120 4.960 74.450 4.975 ;
        RECT 79.445 4.960 79.775 4.975 ;
        RECT 84.780 4.960 85.110 4.975 ;
        RECT 90.105 4.960 90.435 4.975 ;
        RECT 95.440 4.960 95.770 4.975 ;
        RECT 100.765 4.960 101.095 4.975 ;
        RECT 106.100 4.960 106.430 4.975 ;
        RECT 111.425 4.960 111.755 4.975 ;
        RECT 116.760 4.960 117.090 4.975 ;
        RECT 122.085 4.960 122.415 4.975 ;
        RECT 35.980 4.630 36.310 4.645 ;
        RECT 41.305 4.630 41.635 4.645 ;
        RECT 46.640 4.630 46.970 4.645 ;
        RECT 51.965 4.630 52.295 4.645 ;
        RECT 57.300 4.630 57.630 4.645 ;
        RECT 62.625 4.630 62.955 4.645 ;
        RECT 67.960 4.630 68.290 4.645 ;
        RECT 73.285 4.630 73.615 4.645 ;
        RECT 78.620 4.630 78.950 4.645 ;
        RECT 83.945 4.630 84.275 4.645 ;
        RECT 89.280 4.630 89.610 4.645 ;
        RECT 94.605 4.630 94.935 4.645 ;
        RECT 99.940 4.630 100.270 4.645 ;
        RECT 105.265 4.630 105.595 4.645 ;
        RECT 110.600 4.630 110.930 4.645 ;
        RECT 115.925 4.630 116.255 4.645 ;
        RECT 121.260 4.630 121.590 4.645 ;
        RECT 126.585 4.630 126.915 4.645 ;
        RECT 31.240 4.330 127.180 4.630 ;
        RECT 35.980 4.315 36.310 4.330 ;
        RECT 41.305 4.315 41.635 4.330 ;
        RECT 46.640 4.315 46.970 4.330 ;
        RECT 51.965 4.315 52.295 4.330 ;
        RECT 57.300 4.315 57.630 4.330 ;
        RECT 62.625 4.315 62.955 4.330 ;
        RECT 67.960 4.315 68.290 4.330 ;
        RECT 73.285 4.315 73.615 4.330 ;
        RECT 78.620 4.315 78.950 4.330 ;
        RECT 83.945 4.315 84.275 4.330 ;
        RECT 89.280 4.315 89.610 4.330 ;
        RECT 94.605 4.315 94.935 4.330 ;
        RECT 99.940 4.315 100.270 4.330 ;
        RECT 105.265 4.315 105.595 4.330 ;
        RECT 110.600 4.315 110.930 4.330 ;
        RECT 115.925 4.315 116.255 4.330 ;
        RECT 121.260 4.315 121.590 4.330 ;
        RECT 126.585 4.315 126.915 4.330 ;
        RECT 127.670 0.330 129.375 78.415 ;
    END
  END vss
  PIN dvdd
    ANTENNADIFFAREA 7.862400 ;
    PORT
      LAYER nwell ;
        RECT 3.130 60.745 4.665 63.055 ;
        RECT 3.130 52.605 4.665 54.915 ;
        RECT 3.130 44.465 4.665 46.775 ;
        RECT 3.130 36.325 4.665 38.635 ;
        RECT 3.130 28.185 4.665 30.495 ;
        RECT 3.130 20.045 4.665 22.355 ;
        RECT 3.130 11.905 4.665 14.215 ;
        RECT 3.130 3.765 4.665 6.075 ;
      LAYER li1 ;
        RECT 3.675 61.955 4.445 62.930 ;
        RECT 3.765 61.805 4.445 61.955 ;
        RECT 3.765 60.895 4.035 61.805 ;
        RECT 3.675 53.815 4.445 54.790 ;
        RECT 3.765 53.665 4.445 53.815 ;
        RECT 3.765 52.755 4.035 53.665 ;
        RECT 3.675 45.675 4.445 46.650 ;
        RECT 3.765 45.525 4.445 45.675 ;
        RECT 3.765 44.615 4.035 45.525 ;
        RECT 3.675 37.535 4.445 38.510 ;
        RECT 3.765 37.385 4.445 37.535 ;
        RECT 3.765 36.475 4.035 37.385 ;
        RECT 3.675 29.395 4.445 30.370 ;
        RECT 3.765 29.245 4.445 29.395 ;
        RECT 3.765 28.335 4.035 29.245 ;
        RECT 3.675 21.255 4.445 22.230 ;
        RECT 3.765 21.105 4.445 21.255 ;
        RECT 3.765 20.195 4.035 21.105 ;
        RECT 3.675 13.115 4.445 14.090 ;
        RECT 3.765 12.965 4.445 13.115 ;
        RECT 3.765 12.055 4.035 12.965 ;
        RECT 3.675 4.975 4.445 5.950 ;
        RECT 3.765 4.825 4.445 4.975 ;
        RECT 3.765 3.915 4.035 4.825 ;
      LAYER met1 ;
        RECT 0.330 61.750 10.820 62.035 ;
        RECT 0.330 61.535 3.030 61.750 ;
        RECT 0.330 53.610 10.820 53.895 ;
        RECT 0.330 53.395 3.030 53.610 ;
        RECT 0.330 45.470 10.820 45.755 ;
        RECT 0.330 45.255 3.030 45.470 ;
        RECT 0.330 37.330 10.820 37.615 ;
        RECT 0.330 37.115 3.030 37.330 ;
        RECT 0.330 29.190 10.820 29.475 ;
        RECT 0.330 28.975 3.030 29.190 ;
        RECT 0.330 21.050 10.820 21.335 ;
        RECT 0.330 20.835 3.030 21.050 ;
        RECT 0.330 12.910 10.820 13.195 ;
        RECT 0.330 12.695 3.030 12.910 ;
        RECT 0.330 4.770 10.820 5.055 ;
        RECT 0.330 4.555 3.030 4.770 ;
      LAYER met2 ;
        RECT -1.000 71.230 2.985 72.695 ;
        RECT 1.520 1.535 2.985 71.230 ;
    END
  END dvdd
  PIN dvss
    ANTENNADIFFAREA 90.511597 ;
    PORT
      LAYER pwell ;
        RECT 0.200 66.655 22.060 67.085 ;
        RECT 1.955 64.705 6.365 66.655 ;
        RECT 8.755 65.455 10.870 66.655 ;
        RECT 11.040 65.455 14.710 66.655 ;
        RECT 14.995 65.285 21.895 66.655 ;
        RECT 22.825 61.430 24.655 63.260 ;
        RECT 5.420 60.455 9.830 60.895 ;
        RECT 3.185 58.945 9.830 60.455 ;
        RECT 11.160 58.945 13.270 60.190 ;
        RECT 13.555 58.945 20.455 60.315 ;
        RECT 0.200 58.515 22.060 58.945 ;
        RECT 1.955 56.565 6.365 58.515 ;
        RECT 8.755 57.315 10.870 58.515 ;
        RECT 11.040 57.315 14.710 58.515 ;
        RECT 14.995 57.145 21.895 58.515 ;
        RECT 22.825 53.290 24.655 55.120 ;
        RECT 5.420 52.315 9.830 52.755 ;
        RECT 3.185 50.805 9.830 52.315 ;
        RECT 11.160 50.805 13.270 52.050 ;
        RECT 13.555 50.805 20.455 52.175 ;
        RECT 0.200 50.375 22.060 50.805 ;
        RECT 1.955 48.425 6.365 50.375 ;
        RECT 8.755 49.175 10.870 50.375 ;
        RECT 11.040 49.175 14.710 50.375 ;
        RECT 14.995 49.005 21.895 50.375 ;
        RECT 22.825 45.150 24.655 46.980 ;
        RECT 5.420 44.175 9.830 44.615 ;
        RECT 3.185 42.665 9.830 44.175 ;
        RECT 11.160 42.665 13.270 43.910 ;
        RECT 13.555 42.665 20.455 44.035 ;
        RECT 0.200 42.235 22.060 42.665 ;
        RECT 1.955 40.285 6.365 42.235 ;
        RECT 8.755 41.035 10.870 42.235 ;
        RECT 11.040 41.035 14.710 42.235 ;
        RECT 14.995 40.865 21.895 42.235 ;
        RECT 22.825 37.010 24.655 38.840 ;
        RECT 5.420 36.035 9.830 36.475 ;
        RECT 3.185 34.525 9.830 36.035 ;
        RECT 11.160 34.525 13.270 35.770 ;
        RECT 13.555 34.525 20.455 35.895 ;
        RECT 0.200 34.095 22.060 34.525 ;
        RECT 1.955 32.145 6.365 34.095 ;
        RECT 8.755 32.895 10.870 34.095 ;
        RECT 11.040 32.895 14.710 34.095 ;
        RECT 14.995 32.725 21.895 34.095 ;
        RECT 22.825 28.870 24.655 30.700 ;
        RECT 5.420 27.895 9.830 28.335 ;
        RECT 3.185 26.385 9.830 27.895 ;
        RECT 11.160 26.385 13.270 27.630 ;
        RECT 13.555 26.385 20.455 27.755 ;
        RECT 0.200 25.955 22.060 26.385 ;
        RECT 1.955 24.005 6.365 25.955 ;
        RECT 8.755 24.755 10.870 25.955 ;
        RECT 11.040 24.755 14.710 25.955 ;
        RECT 14.995 24.585 21.895 25.955 ;
        RECT 22.825 20.730 24.655 22.560 ;
        RECT 5.420 19.755 9.830 20.195 ;
        RECT 3.185 18.245 9.830 19.755 ;
        RECT 11.160 18.245 13.270 19.490 ;
        RECT 13.555 18.245 20.455 19.615 ;
        RECT 0.200 17.815 22.060 18.245 ;
        RECT 1.955 15.865 6.365 17.815 ;
        RECT 8.755 16.615 10.870 17.815 ;
        RECT 11.040 16.615 14.710 17.815 ;
        RECT 14.995 16.445 21.895 17.815 ;
        RECT 22.825 12.590 24.655 14.420 ;
        RECT 5.420 11.615 9.830 12.055 ;
        RECT 3.185 10.105 9.830 11.615 ;
        RECT 11.160 10.105 13.270 11.350 ;
        RECT 13.555 10.105 20.455 11.475 ;
        RECT 0.200 9.675 22.060 10.105 ;
        RECT 1.955 7.725 6.365 9.675 ;
        RECT 8.755 8.475 10.870 9.675 ;
        RECT 11.040 8.475 14.710 9.675 ;
        RECT 14.995 8.305 21.895 9.675 ;
        RECT 22.825 4.450 24.655 6.280 ;
        RECT 5.420 3.475 9.830 3.915 ;
        RECT 3.185 1.965 9.830 3.475 ;
        RECT 11.160 1.965 13.270 3.210 ;
        RECT 13.555 1.965 20.455 3.335 ;
        RECT 0.200 1.535 22.060 1.965 ;
      LAYER li1 ;
        RECT 0.330 66.785 21.930 66.955 ;
        RECT 1.915 66.445 5.625 66.615 ;
        RECT 1.915 64.815 2.505 66.445 ;
        RECT 3.475 64.895 4.065 66.445 ;
        RECT 5.035 64.895 5.625 66.445 ;
        RECT 9.540 65.565 10.130 66.475 ;
        RECT 10.980 65.545 11.570 66.505 ;
        RECT 12.360 65.820 13.310 66.505 ;
        RECT 14.270 65.545 14.600 66.505 ;
        RECT 14.825 66.320 21.835 66.490 ;
        RECT 14.825 65.485 15.715 66.320 ;
        RECT 16.305 65.825 17.315 66.320 ;
        RECT 17.865 65.825 18.875 66.320 ;
        RECT 19.425 65.825 20.475 66.320 ;
        RECT 21.465 65.825 21.835 66.320 ;
        RECT 23.005 62.910 24.475 63.080 ;
        RECT 23.005 61.780 23.175 62.910 ;
        RECT 24.305 61.780 24.475 62.910 ;
        RECT 23.005 61.610 24.475 61.780 ;
        RECT 3.765 59.295 4.035 60.305 ;
        RECT 3.425 59.065 4.375 59.295 ;
        RECT 5.380 59.155 5.970 60.705 ;
        RECT 6.940 59.155 7.530 60.705 ;
        RECT 8.500 59.155 9.090 60.705 ;
        RECT 5.380 58.985 9.090 59.155 ;
        RECT 10.980 59.095 11.910 60.100 ;
        RECT 12.870 59.095 13.200 60.100 ;
        RECT 13.385 59.280 14.275 60.115 ;
        RECT 14.865 59.280 15.875 59.775 ;
        RECT 16.425 59.280 17.435 59.775 ;
        RECT 17.985 59.280 19.035 59.775 ;
        RECT 20.025 59.280 20.395 59.775 ;
        RECT 13.385 59.110 20.395 59.280 ;
        RECT 0.330 58.645 21.930 58.815 ;
        RECT 1.915 58.305 5.625 58.475 ;
        RECT 1.915 56.675 2.505 58.305 ;
        RECT 3.475 56.755 4.065 58.305 ;
        RECT 5.035 56.755 5.625 58.305 ;
        RECT 9.540 57.425 10.130 58.335 ;
        RECT 10.980 57.405 11.570 58.365 ;
        RECT 12.360 57.680 13.310 58.365 ;
        RECT 14.270 57.405 14.600 58.365 ;
        RECT 14.825 58.180 21.835 58.350 ;
        RECT 14.825 57.345 15.715 58.180 ;
        RECT 16.305 57.685 17.315 58.180 ;
        RECT 17.865 57.685 18.875 58.180 ;
        RECT 19.425 57.685 20.475 58.180 ;
        RECT 21.465 57.685 21.835 58.180 ;
        RECT 23.005 54.770 24.475 54.940 ;
        RECT 23.005 53.640 23.175 54.770 ;
        RECT 24.305 53.640 24.475 54.770 ;
        RECT 23.005 53.470 24.475 53.640 ;
        RECT 3.765 51.155 4.035 52.165 ;
        RECT 3.425 50.925 4.375 51.155 ;
        RECT 5.380 51.015 5.970 52.565 ;
        RECT 6.940 51.015 7.530 52.565 ;
        RECT 8.500 51.015 9.090 52.565 ;
        RECT 5.380 50.845 9.090 51.015 ;
        RECT 10.980 50.955 11.910 51.960 ;
        RECT 12.870 50.955 13.200 51.960 ;
        RECT 13.385 51.140 14.275 51.975 ;
        RECT 14.865 51.140 15.875 51.635 ;
        RECT 16.425 51.140 17.435 51.635 ;
        RECT 17.985 51.140 19.035 51.635 ;
        RECT 20.025 51.140 20.395 51.635 ;
        RECT 13.385 50.970 20.395 51.140 ;
        RECT 0.330 50.505 21.930 50.675 ;
        RECT 1.915 50.165 5.625 50.335 ;
        RECT 1.915 48.535 2.505 50.165 ;
        RECT 3.475 48.615 4.065 50.165 ;
        RECT 5.035 48.615 5.625 50.165 ;
        RECT 9.540 49.285 10.130 50.195 ;
        RECT 10.980 49.265 11.570 50.225 ;
        RECT 12.360 49.540 13.310 50.225 ;
        RECT 14.270 49.265 14.600 50.225 ;
        RECT 14.825 50.040 21.835 50.210 ;
        RECT 14.825 49.205 15.715 50.040 ;
        RECT 16.305 49.545 17.315 50.040 ;
        RECT 17.865 49.545 18.875 50.040 ;
        RECT 19.425 49.545 20.475 50.040 ;
        RECT 21.465 49.545 21.835 50.040 ;
        RECT 23.005 46.630 24.475 46.800 ;
        RECT 23.005 45.500 23.175 46.630 ;
        RECT 24.305 45.500 24.475 46.630 ;
        RECT 23.005 45.330 24.475 45.500 ;
        RECT 3.765 43.015 4.035 44.025 ;
        RECT 3.425 42.785 4.375 43.015 ;
        RECT 5.380 42.875 5.970 44.425 ;
        RECT 6.940 42.875 7.530 44.425 ;
        RECT 8.500 42.875 9.090 44.425 ;
        RECT 5.380 42.705 9.090 42.875 ;
        RECT 10.980 42.815 11.910 43.820 ;
        RECT 12.870 42.815 13.200 43.820 ;
        RECT 13.385 43.000 14.275 43.835 ;
        RECT 14.865 43.000 15.875 43.495 ;
        RECT 16.425 43.000 17.435 43.495 ;
        RECT 17.985 43.000 19.035 43.495 ;
        RECT 20.025 43.000 20.395 43.495 ;
        RECT 13.385 42.830 20.395 43.000 ;
        RECT 0.330 42.365 21.930 42.535 ;
        RECT 1.915 42.025 5.625 42.195 ;
        RECT 1.915 40.395 2.505 42.025 ;
        RECT 3.475 40.475 4.065 42.025 ;
        RECT 5.035 40.475 5.625 42.025 ;
        RECT 9.540 41.145 10.130 42.055 ;
        RECT 10.980 41.125 11.570 42.085 ;
        RECT 12.360 41.400 13.310 42.085 ;
        RECT 14.270 41.125 14.600 42.085 ;
        RECT 14.825 41.900 21.835 42.070 ;
        RECT 14.825 41.065 15.715 41.900 ;
        RECT 16.305 41.405 17.315 41.900 ;
        RECT 17.865 41.405 18.875 41.900 ;
        RECT 19.425 41.405 20.475 41.900 ;
        RECT 21.465 41.405 21.835 41.900 ;
        RECT 23.005 38.490 24.475 38.660 ;
        RECT 23.005 37.360 23.175 38.490 ;
        RECT 24.305 37.360 24.475 38.490 ;
        RECT 23.005 37.190 24.475 37.360 ;
        RECT 3.765 34.875 4.035 35.885 ;
        RECT 3.425 34.645 4.375 34.875 ;
        RECT 5.380 34.735 5.970 36.285 ;
        RECT 6.940 34.735 7.530 36.285 ;
        RECT 8.500 34.735 9.090 36.285 ;
        RECT 5.380 34.565 9.090 34.735 ;
        RECT 10.980 34.675 11.910 35.680 ;
        RECT 12.870 34.675 13.200 35.680 ;
        RECT 13.385 34.860 14.275 35.695 ;
        RECT 14.865 34.860 15.875 35.355 ;
        RECT 16.425 34.860 17.435 35.355 ;
        RECT 17.985 34.860 19.035 35.355 ;
        RECT 20.025 34.860 20.395 35.355 ;
        RECT 13.385 34.690 20.395 34.860 ;
        RECT 0.330 34.225 21.930 34.395 ;
        RECT 1.915 33.885 5.625 34.055 ;
        RECT 1.915 32.255 2.505 33.885 ;
        RECT 3.475 32.335 4.065 33.885 ;
        RECT 5.035 32.335 5.625 33.885 ;
        RECT 9.540 33.005 10.130 33.915 ;
        RECT 10.980 32.985 11.570 33.945 ;
        RECT 12.360 33.260 13.310 33.945 ;
        RECT 14.270 32.985 14.600 33.945 ;
        RECT 14.825 33.760 21.835 33.930 ;
        RECT 14.825 32.925 15.715 33.760 ;
        RECT 16.305 33.265 17.315 33.760 ;
        RECT 17.865 33.265 18.875 33.760 ;
        RECT 19.425 33.265 20.475 33.760 ;
        RECT 21.465 33.265 21.835 33.760 ;
        RECT 23.005 30.350 24.475 30.520 ;
        RECT 23.005 29.220 23.175 30.350 ;
        RECT 24.305 29.220 24.475 30.350 ;
        RECT 23.005 29.050 24.475 29.220 ;
        RECT 3.765 26.735 4.035 27.745 ;
        RECT 3.425 26.505 4.375 26.735 ;
        RECT 5.380 26.595 5.970 28.145 ;
        RECT 6.940 26.595 7.530 28.145 ;
        RECT 8.500 26.595 9.090 28.145 ;
        RECT 5.380 26.425 9.090 26.595 ;
        RECT 10.980 26.535 11.910 27.540 ;
        RECT 12.870 26.535 13.200 27.540 ;
        RECT 13.385 26.720 14.275 27.555 ;
        RECT 14.865 26.720 15.875 27.215 ;
        RECT 16.425 26.720 17.435 27.215 ;
        RECT 17.985 26.720 19.035 27.215 ;
        RECT 20.025 26.720 20.395 27.215 ;
        RECT 13.385 26.550 20.395 26.720 ;
        RECT 0.330 26.085 21.930 26.255 ;
        RECT 1.915 25.745 5.625 25.915 ;
        RECT 1.915 24.115 2.505 25.745 ;
        RECT 3.475 24.195 4.065 25.745 ;
        RECT 5.035 24.195 5.625 25.745 ;
        RECT 9.540 24.865 10.130 25.775 ;
        RECT 10.980 24.845 11.570 25.805 ;
        RECT 12.360 25.120 13.310 25.805 ;
        RECT 14.270 24.845 14.600 25.805 ;
        RECT 14.825 25.620 21.835 25.790 ;
        RECT 14.825 24.785 15.715 25.620 ;
        RECT 16.305 25.125 17.315 25.620 ;
        RECT 17.865 25.125 18.875 25.620 ;
        RECT 19.425 25.125 20.475 25.620 ;
        RECT 21.465 25.125 21.835 25.620 ;
        RECT 23.005 22.210 24.475 22.380 ;
        RECT 23.005 21.080 23.175 22.210 ;
        RECT 24.305 21.080 24.475 22.210 ;
        RECT 23.005 20.910 24.475 21.080 ;
        RECT 3.765 18.595 4.035 19.605 ;
        RECT 3.425 18.365 4.375 18.595 ;
        RECT 5.380 18.455 5.970 20.005 ;
        RECT 6.940 18.455 7.530 20.005 ;
        RECT 8.500 18.455 9.090 20.005 ;
        RECT 5.380 18.285 9.090 18.455 ;
        RECT 10.980 18.395 11.910 19.400 ;
        RECT 12.870 18.395 13.200 19.400 ;
        RECT 13.385 18.580 14.275 19.415 ;
        RECT 14.865 18.580 15.875 19.075 ;
        RECT 16.425 18.580 17.435 19.075 ;
        RECT 17.985 18.580 19.035 19.075 ;
        RECT 20.025 18.580 20.395 19.075 ;
        RECT 13.385 18.410 20.395 18.580 ;
        RECT 0.330 17.945 21.930 18.115 ;
        RECT 1.915 17.605 5.625 17.775 ;
        RECT 1.915 15.975 2.505 17.605 ;
        RECT 3.475 16.055 4.065 17.605 ;
        RECT 5.035 16.055 5.625 17.605 ;
        RECT 9.540 16.725 10.130 17.635 ;
        RECT 10.980 16.705 11.570 17.665 ;
        RECT 12.360 16.980 13.310 17.665 ;
        RECT 14.270 16.705 14.600 17.665 ;
        RECT 14.825 17.480 21.835 17.650 ;
        RECT 14.825 16.645 15.715 17.480 ;
        RECT 16.305 16.985 17.315 17.480 ;
        RECT 17.865 16.985 18.875 17.480 ;
        RECT 19.425 16.985 20.475 17.480 ;
        RECT 21.465 16.985 21.835 17.480 ;
        RECT 23.005 14.070 24.475 14.240 ;
        RECT 23.005 12.940 23.175 14.070 ;
        RECT 24.305 12.940 24.475 14.070 ;
        RECT 23.005 12.770 24.475 12.940 ;
        RECT 3.765 10.455 4.035 11.465 ;
        RECT 3.425 10.225 4.375 10.455 ;
        RECT 5.380 10.315 5.970 11.865 ;
        RECT 6.940 10.315 7.530 11.865 ;
        RECT 8.500 10.315 9.090 11.865 ;
        RECT 5.380 10.145 9.090 10.315 ;
        RECT 10.980 10.255 11.910 11.260 ;
        RECT 12.870 10.255 13.200 11.260 ;
        RECT 13.385 10.440 14.275 11.275 ;
        RECT 14.865 10.440 15.875 10.935 ;
        RECT 16.425 10.440 17.435 10.935 ;
        RECT 17.985 10.440 19.035 10.935 ;
        RECT 20.025 10.440 20.395 10.935 ;
        RECT 13.385 10.270 20.395 10.440 ;
        RECT 0.330 9.805 21.930 9.975 ;
        RECT 1.915 9.465 5.625 9.635 ;
        RECT 1.915 7.835 2.505 9.465 ;
        RECT 3.475 7.915 4.065 9.465 ;
        RECT 5.035 7.915 5.625 9.465 ;
        RECT 9.540 8.585 10.130 9.495 ;
        RECT 10.980 8.565 11.570 9.525 ;
        RECT 12.360 8.840 13.310 9.525 ;
        RECT 14.270 8.565 14.600 9.525 ;
        RECT 14.825 9.340 21.835 9.510 ;
        RECT 14.825 8.505 15.715 9.340 ;
        RECT 16.305 8.845 17.315 9.340 ;
        RECT 17.865 8.845 18.875 9.340 ;
        RECT 19.425 8.845 20.475 9.340 ;
        RECT 21.465 8.845 21.835 9.340 ;
        RECT 23.005 5.930 24.475 6.100 ;
        RECT 23.005 4.800 23.175 5.930 ;
        RECT 24.305 4.800 24.475 5.930 ;
        RECT 23.005 4.630 24.475 4.800 ;
        RECT 3.765 2.315 4.035 3.325 ;
        RECT 3.425 2.085 4.375 2.315 ;
        RECT 5.380 2.175 5.970 3.725 ;
        RECT 6.940 2.175 7.530 3.725 ;
        RECT 8.500 2.175 9.090 3.725 ;
        RECT 5.380 2.005 9.090 2.175 ;
        RECT 10.980 2.115 11.910 3.120 ;
        RECT 12.870 2.115 13.200 3.120 ;
        RECT 13.385 2.300 14.275 3.135 ;
        RECT 14.865 2.300 15.875 2.795 ;
        RECT 16.425 2.300 17.435 2.795 ;
        RECT 17.985 2.300 19.035 2.795 ;
        RECT 20.025 2.300 20.395 2.795 ;
        RECT 13.385 2.130 20.395 2.300 ;
        RECT 0.330 1.665 21.930 1.835 ;
      LAYER met1 ;
        RECT 0.330 66.245 21.930 66.985 ;
        RECT 23.340 62.790 24.510 63.110 ;
        RECT 24.160 61.510 24.510 62.790 ;
        RECT 13.910 61.190 24.510 61.510 ;
        RECT 13.910 59.355 14.235 61.190 ;
        RECT 0.330 58.105 21.930 59.355 ;
        RECT 23.340 54.650 24.510 54.970 ;
        RECT 24.160 53.370 24.510 54.650 ;
        RECT 13.910 53.050 24.510 53.370 ;
        RECT 13.910 51.215 14.235 53.050 ;
        RECT 0.330 49.965 21.930 51.215 ;
        RECT 23.340 46.510 24.510 46.830 ;
        RECT 24.160 45.230 24.510 46.510 ;
        RECT 13.910 44.910 24.510 45.230 ;
        RECT 13.910 43.075 14.235 44.910 ;
        RECT 0.330 41.825 21.930 43.075 ;
        RECT 23.340 38.370 24.510 38.690 ;
        RECT 24.160 37.090 24.510 38.370 ;
        RECT 13.910 36.770 24.510 37.090 ;
        RECT 13.910 34.935 14.235 36.770 ;
        RECT 0.330 33.685 21.930 34.935 ;
        RECT 23.340 30.230 24.510 30.550 ;
        RECT 24.160 28.950 24.510 30.230 ;
        RECT 13.910 28.630 24.510 28.950 ;
        RECT 13.910 26.795 14.235 28.630 ;
        RECT 0.330 25.545 21.930 26.795 ;
        RECT 23.340 22.090 24.510 22.410 ;
        RECT 24.160 20.810 24.510 22.090 ;
        RECT 13.910 20.490 24.510 20.810 ;
        RECT 13.910 18.655 14.235 20.490 ;
        RECT 0.330 17.405 21.930 18.655 ;
        RECT 23.340 13.950 24.510 14.270 ;
        RECT 24.160 12.670 24.510 13.950 ;
        RECT 13.910 12.350 24.510 12.670 ;
        RECT 13.910 10.515 14.235 12.350 ;
        RECT 0.330 9.265 21.930 10.515 ;
        RECT 23.340 5.810 24.510 6.130 ;
        RECT 24.160 4.530 24.510 5.810 ;
        RECT 13.910 4.210 24.510 4.530 ;
        RECT 13.910 2.375 14.235 4.210 ;
        RECT 0.330 1.635 21.930 2.375 ;
      LAYER met2 ;
        RECT -1.000 73.455 9.055 75.350 ;
        RECT 7.160 1.510 9.055 73.455 ;
    END
  END dvss
  PIN Vhigh
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER li1 ;
        RECT 38.050 12.070 38.220 12.760 ;
        RECT 34.895 7.720 35.065 8.760 ;
        RECT 35.610 7.280 36.320 11.855 ;
        RECT 36.800 7.265 37.510 11.840 ;
        RECT 38.050 10.275 38.220 11.315 ;
        RECT 34.895 6.275 35.065 6.965 ;
      LAYER met1 ;
        RECT 36.020 10.235 36.375 11.855 ;
        RECT 36.745 10.235 37.100 11.840 ;
        RECT 38.020 11.775 38.250 12.740 ;
        RECT 36.020 9.645 37.100 10.235 ;
        RECT 37.240 11.605 38.250 11.775 ;
        RECT 37.240 9.645 37.410 11.605 ;
        RECT 38.020 10.295 38.250 11.605 ;
        RECT 35.705 9.370 37.410 9.645 ;
        RECT 34.865 7.430 35.095 8.740 ;
        RECT 35.705 7.430 35.875 9.370 ;
        RECT 34.865 7.260 35.875 7.430 ;
        RECT 36.020 7.265 37.100 9.370 ;
        RECT 34.865 6.295 35.095 7.260 ;
        RECT 36.020 7.215 37.095 7.265 ;
      LAYER met2 ;
        RECT 34.685 7.215 37.095 7.650 ;
      LAYER met3 ;
        RECT 34.480 -0.020 35.665 7.675 ;
    END
  END Vhigh
  PIN Vlow
    ANTENNADIFFAREA 0.957000 ;
    PORT
      LAYER li1 ;
        RECT 123.330 12.070 123.500 12.760 ;
        RECT 120.175 7.720 120.345 8.760 ;
        RECT 120.890 7.260 121.600 11.835 ;
        RECT 122.080 7.280 122.790 11.855 ;
        RECT 123.330 10.275 123.500 11.315 ;
        RECT 120.175 6.275 120.345 6.965 ;
      LAYER met1 ;
        RECT 121.300 10.235 121.655 11.835 ;
        RECT 121.300 10.230 121.845 10.235 ;
        RECT 122.025 10.230 122.380 11.855 ;
        RECT 123.300 11.775 123.530 12.740 ;
        RECT 121.300 9.645 122.380 10.230 ;
        RECT 122.520 11.605 123.530 11.775 ;
        RECT 122.520 9.645 122.690 11.605 ;
        RECT 123.300 10.295 123.530 11.605 ;
        RECT 120.985 9.370 122.690 9.645 ;
        RECT 120.145 7.430 120.375 8.740 ;
        RECT 120.985 7.430 121.155 9.370 ;
        RECT 120.145 7.260 121.155 7.430 ;
        RECT 121.300 7.280 122.380 9.370 ;
        RECT 120.145 6.295 120.375 7.260 ;
        RECT 121.300 7.215 122.375 7.280 ;
      LAYER met2 ;
        RECT 122.510 7.715 123.510 8.150 ;
        RECT 122.510 7.650 122.945 7.715 ;
        RECT 121.300 7.215 122.945 7.650 ;
      LAYER met3 ;
        RECT 122.735 -0.020 123.840 8.175 ;
    END
  END Vlow
  OBS
      LAYER li1 ;
        RECT 31.475 75.095 32.185 77.380 ;
        RECT 32.725 75.535 32.895 76.575 ;
        RECT 33.515 75.535 33.685 76.575 ;
        RECT 34.105 75.535 34.275 76.575 ;
        RECT 34.895 75.535 35.065 76.575 ;
        RECT 35.610 75.095 36.320 77.380 ;
        RECT 36.800 75.080 37.510 77.365 ;
        RECT 38.050 75.535 38.220 76.575 ;
        RECT 38.840 75.535 39.010 76.575 ;
        RECT 39.430 75.535 39.600 76.575 ;
        RECT 40.220 75.535 40.390 76.575 ;
        RECT 40.935 75.075 41.645 77.360 ;
        RECT 42.135 75.080 42.845 77.365 ;
        RECT 43.385 75.535 43.555 76.575 ;
        RECT 44.175 75.535 44.345 76.575 ;
        RECT 44.765 75.535 44.935 76.575 ;
        RECT 45.555 75.535 45.725 76.575 ;
        RECT 46.270 75.075 46.980 77.360 ;
        RECT 47.460 75.080 48.170 77.365 ;
        RECT 48.710 75.535 48.880 76.575 ;
        RECT 49.500 75.535 49.670 76.575 ;
        RECT 50.090 75.535 50.260 76.575 ;
        RECT 50.880 75.535 51.050 76.575 ;
        RECT 51.595 75.075 52.305 77.360 ;
        RECT 52.795 75.080 53.505 77.365 ;
        RECT 54.045 75.535 54.215 76.575 ;
        RECT 54.835 75.535 55.005 76.575 ;
        RECT 55.425 75.535 55.595 76.575 ;
        RECT 56.215 75.535 56.385 76.575 ;
        RECT 56.930 75.075 57.640 77.360 ;
        RECT 58.120 75.080 58.830 77.365 ;
        RECT 59.370 75.535 59.540 76.575 ;
        RECT 60.160 75.535 60.330 76.575 ;
        RECT 60.750 75.535 60.920 76.575 ;
        RECT 61.540 75.535 61.710 76.575 ;
        RECT 62.255 75.075 62.965 77.360 ;
        RECT 63.455 75.080 64.165 77.365 ;
        RECT 64.705 75.535 64.875 76.575 ;
        RECT 65.495 75.535 65.665 76.575 ;
        RECT 66.085 75.535 66.255 76.575 ;
        RECT 66.875 75.535 67.045 76.575 ;
        RECT 67.590 75.075 68.300 77.360 ;
        RECT 68.780 75.080 69.490 77.365 ;
        RECT 70.030 75.535 70.200 76.575 ;
        RECT 70.820 75.535 70.990 76.575 ;
        RECT 71.410 75.535 71.580 76.575 ;
        RECT 72.200 75.535 72.370 76.575 ;
        RECT 72.915 75.075 73.625 77.360 ;
        RECT 74.115 75.080 74.825 77.365 ;
        RECT 75.365 75.535 75.535 76.575 ;
        RECT 76.155 75.535 76.325 76.575 ;
        RECT 76.745 75.535 76.915 76.575 ;
        RECT 77.535 75.535 77.705 76.575 ;
        RECT 78.250 75.075 78.960 77.360 ;
        RECT 79.440 75.080 80.150 77.365 ;
        RECT 80.690 75.535 80.860 76.575 ;
        RECT 81.480 75.535 81.650 76.575 ;
        RECT 82.070 75.535 82.240 76.575 ;
        RECT 82.860 75.535 83.030 76.575 ;
        RECT 83.575 75.075 84.285 77.360 ;
        RECT 84.775 75.080 85.485 77.365 ;
        RECT 86.025 75.535 86.195 76.575 ;
        RECT 86.815 75.535 86.985 76.575 ;
        RECT 87.405 75.535 87.575 76.575 ;
        RECT 88.195 75.535 88.365 76.575 ;
        RECT 88.910 75.075 89.620 77.360 ;
        RECT 90.100 75.080 90.810 77.365 ;
        RECT 91.350 75.535 91.520 76.575 ;
        RECT 92.140 75.535 92.310 76.575 ;
        RECT 92.730 75.535 92.900 76.575 ;
        RECT 93.520 75.535 93.690 76.575 ;
        RECT 94.235 75.075 94.945 77.360 ;
        RECT 95.435 75.080 96.145 77.365 ;
        RECT 96.685 75.535 96.855 76.575 ;
        RECT 97.475 75.535 97.645 76.575 ;
        RECT 98.065 75.535 98.235 76.575 ;
        RECT 98.855 75.535 99.025 76.575 ;
        RECT 99.570 75.075 100.280 77.360 ;
        RECT 100.760 75.080 101.470 77.365 ;
        RECT 102.010 75.535 102.180 76.575 ;
        RECT 102.800 75.535 102.970 76.575 ;
        RECT 103.390 75.535 103.560 76.575 ;
        RECT 104.180 75.535 104.350 76.575 ;
        RECT 104.895 75.075 105.605 77.360 ;
        RECT 106.095 75.080 106.805 77.365 ;
        RECT 107.345 75.535 107.515 76.575 ;
        RECT 108.135 75.535 108.305 76.575 ;
        RECT 108.725 75.535 108.895 76.575 ;
        RECT 109.515 75.535 109.685 76.575 ;
        RECT 110.230 75.075 110.940 77.360 ;
        RECT 111.420 75.080 112.130 77.365 ;
        RECT 112.670 75.535 112.840 76.575 ;
        RECT 113.460 75.535 113.630 76.575 ;
        RECT 114.050 75.535 114.220 76.575 ;
        RECT 114.840 75.535 115.010 76.575 ;
        RECT 115.555 75.075 116.265 77.360 ;
        RECT 116.755 75.080 117.465 77.365 ;
        RECT 118.005 75.535 118.175 76.575 ;
        RECT 118.795 75.535 118.965 76.575 ;
        RECT 119.385 75.535 119.555 76.575 ;
        RECT 120.175 75.535 120.345 76.575 ;
        RECT 120.890 75.075 121.600 77.360 ;
        RECT 122.080 75.095 122.790 77.380 ;
        RECT 123.330 75.535 123.500 76.575 ;
        RECT 124.120 75.535 124.290 76.575 ;
        RECT 124.710 75.535 124.880 76.575 ;
        RECT 125.500 75.535 125.670 76.575 ;
        RECT 126.215 75.095 126.925 77.380 ;
        RECT 32.725 74.090 32.895 74.780 ;
        RECT 33.515 74.090 33.685 74.780 ;
        RECT 34.105 74.090 34.275 74.780 ;
        RECT 34.895 74.090 35.065 74.780 ;
        RECT 38.050 74.090 38.220 74.780 ;
        RECT 38.840 74.090 39.010 74.780 ;
        RECT 39.430 74.090 39.600 74.780 ;
        RECT 40.220 74.090 40.390 74.780 ;
        RECT 43.385 74.090 43.555 74.780 ;
        RECT 44.175 74.090 44.345 74.780 ;
        RECT 44.765 74.090 44.935 74.780 ;
        RECT 45.555 74.090 45.725 74.780 ;
        RECT 48.710 74.090 48.880 74.780 ;
        RECT 49.500 74.090 49.670 74.780 ;
        RECT 50.090 74.090 50.260 74.780 ;
        RECT 50.880 74.090 51.050 74.780 ;
        RECT 54.045 74.090 54.215 74.780 ;
        RECT 54.835 74.090 55.005 74.780 ;
        RECT 55.425 74.090 55.595 74.780 ;
        RECT 56.215 74.090 56.385 74.780 ;
        RECT 59.370 74.090 59.540 74.780 ;
        RECT 60.160 74.090 60.330 74.780 ;
        RECT 60.750 74.090 60.920 74.780 ;
        RECT 61.540 74.090 61.710 74.780 ;
        RECT 64.705 74.090 64.875 74.780 ;
        RECT 65.495 74.090 65.665 74.780 ;
        RECT 66.085 74.090 66.255 74.780 ;
        RECT 66.875 74.090 67.045 74.780 ;
        RECT 70.030 74.090 70.200 74.780 ;
        RECT 70.820 74.090 70.990 74.780 ;
        RECT 71.410 74.090 71.580 74.780 ;
        RECT 72.200 74.090 72.370 74.780 ;
        RECT 75.365 74.090 75.535 74.780 ;
        RECT 76.155 74.090 76.325 74.780 ;
        RECT 76.745 74.090 76.915 74.780 ;
        RECT 77.535 74.090 77.705 74.780 ;
        RECT 80.690 74.090 80.860 74.780 ;
        RECT 81.480 74.090 81.650 74.780 ;
        RECT 82.070 74.090 82.240 74.780 ;
        RECT 82.860 74.090 83.030 74.780 ;
        RECT 86.025 74.090 86.195 74.780 ;
        RECT 86.815 74.090 86.985 74.780 ;
        RECT 87.405 74.090 87.575 74.780 ;
        RECT 88.195 74.090 88.365 74.780 ;
        RECT 91.350 74.090 91.520 74.780 ;
        RECT 92.140 74.090 92.310 74.780 ;
        RECT 92.730 74.090 92.900 74.780 ;
        RECT 93.520 74.090 93.690 74.780 ;
        RECT 96.685 74.090 96.855 74.780 ;
        RECT 97.475 74.090 97.645 74.780 ;
        RECT 98.065 74.090 98.235 74.780 ;
        RECT 98.855 74.090 99.025 74.780 ;
        RECT 102.010 74.090 102.180 74.780 ;
        RECT 102.800 74.090 102.970 74.780 ;
        RECT 103.390 74.090 103.560 74.780 ;
        RECT 104.180 74.090 104.350 74.780 ;
        RECT 107.345 74.090 107.515 74.780 ;
        RECT 108.135 74.090 108.305 74.780 ;
        RECT 108.725 74.090 108.895 74.780 ;
        RECT 109.515 74.090 109.685 74.780 ;
        RECT 112.670 74.090 112.840 74.780 ;
        RECT 113.460 74.090 113.630 74.780 ;
        RECT 114.050 74.090 114.220 74.780 ;
        RECT 114.840 74.090 115.010 74.780 ;
        RECT 118.005 74.090 118.175 74.780 ;
        RECT 118.795 74.090 118.965 74.780 ;
        RECT 119.385 74.090 119.555 74.780 ;
        RECT 120.175 74.090 120.345 74.780 ;
        RECT 123.330 74.090 123.500 74.780 ;
        RECT 124.120 74.090 124.290 74.780 ;
        RECT 124.710 74.090 124.880 74.780 ;
        RECT 125.500 74.090 125.670 74.780 ;
        RECT 32.725 72.350 32.895 73.040 ;
        RECT 33.515 72.350 33.685 73.040 ;
        RECT 34.105 72.350 34.275 73.040 ;
        RECT 34.895 72.350 35.065 73.040 ;
        RECT 38.050 72.350 38.220 73.040 ;
        RECT 38.840 72.350 39.010 73.040 ;
        RECT 39.430 72.350 39.600 73.040 ;
        RECT 40.220 72.350 40.390 73.040 ;
        RECT 43.385 72.350 43.555 73.040 ;
        RECT 44.175 72.350 44.345 73.040 ;
        RECT 44.765 72.350 44.935 73.040 ;
        RECT 45.555 72.350 45.725 73.040 ;
        RECT 48.710 72.350 48.880 73.040 ;
        RECT 49.500 72.350 49.670 73.040 ;
        RECT 50.090 72.350 50.260 73.040 ;
        RECT 50.880 72.350 51.050 73.040 ;
        RECT 54.045 72.350 54.215 73.040 ;
        RECT 54.835 72.350 55.005 73.040 ;
        RECT 55.425 72.350 55.595 73.040 ;
        RECT 56.215 72.350 56.385 73.040 ;
        RECT 59.370 72.350 59.540 73.040 ;
        RECT 60.160 72.350 60.330 73.040 ;
        RECT 60.750 72.350 60.920 73.040 ;
        RECT 61.540 72.350 61.710 73.040 ;
        RECT 64.705 72.350 64.875 73.040 ;
        RECT 65.495 72.350 65.665 73.040 ;
        RECT 66.085 72.350 66.255 73.040 ;
        RECT 66.875 72.350 67.045 73.040 ;
        RECT 70.030 72.350 70.200 73.040 ;
        RECT 70.820 72.350 70.990 73.040 ;
        RECT 71.410 72.350 71.580 73.040 ;
        RECT 72.200 72.350 72.370 73.040 ;
        RECT 75.365 72.350 75.535 73.040 ;
        RECT 76.155 72.350 76.325 73.040 ;
        RECT 76.745 72.350 76.915 73.040 ;
        RECT 77.535 72.350 77.705 73.040 ;
        RECT 80.690 72.350 80.860 73.040 ;
        RECT 81.480 72.350 81.650 73.040 ;
        RECT 82.070 72.350 82.240 73.040 ;
        RECT 82.860 72.350 83.030 73.040 ;
        RECT 86.025 72.350 86.195 73.040 ;
        RECT 86.815 72.350 86.985 73.040 ;
        RECT 87.405 72.350 87.575 73.040 ;
        RECT 88.195 72.350 88.365 73.040 ;
        RECT 91.350 72.350 91.520 73.040 ;
        RECT 92.140 72.350 92.310 73.040 ;
        RECT 92.730 72.350 92.900 73.040 ;
        RECT 93.520 72.350 93.690 73.040 ;
        RECT 96.685 72.350 96.855 73.040 ;
        RECT 97.475 72.350 97.645 73.040 ;
        RECT 98.065 72.350 98.235 73.040 ;
        RECT 98.855 72.350 99.025 73.040 ;
        RECT 102.010 72.350 102.180 73.040 ;
        RECT 102.800 72.350 102.970 73.040 ;
        RECT 103.390 72.350 103.560 73.040 ;
        RECT 104.180 72.350 104.350 73.040 ;
        RECT 107.345 72.350 107.515 73.040 ;
        RECT 108.135 72.350 108.305 73.040 ;
        RECT 108.725 72.350 108.895 73.040 ;
        RECT 109.515 72.350 109.685 73.040 ;
        RECT 112.670 72.350 112.840 73.040 ;
        RECT 113.460 72.350 113.630 73.040 ;
        RECT 114.050 72.350 114.220 73.040 ;
        RECT 114.840 72.350 115.010 73.040 ;
        RECT 118.005 72.350 118.175 73.040 ;
        RECT 118.795 72.350 118.965 73.040 ;
        RECT 119.385 72.350 119.555 73.040 ;
        RECT 120.175 72.350 120.345 73.040 ;
        RECT 123.330 72.350 123.500 73.040 ;
        RECT 124.120 72.350 124.290 73.040 ;
        RECT 124.710 72.350 124.880 73.040 ;
        RECT 125.500 72.350 125.670 73.040 ;
        RECT 31.475 67.560 32.185 72.135 ;
        RECT 32.725 70.555 32.895 71.595 ;
        RECT 33.515 70.555 33.685 71.595 ;
        RECT 34.105 70.555 34.275 71.595 ;
        RECT 34.895 70.555 35.065 71.595 ;
        RECT 32.725 68.000 32.895 69.040 ;
        RECT 33.515 68.000 33.685 69.040 ;
        RECT 34.105 68.000 34.275 69.040 ;
        RECT 34.895 68.000 35.065 69.040 ;
        RECT 35.610 67.560 36.320 72.135 ;
        RECT 36.800 67.545 37.510 72.120 ;
        RECT 38.050 70.555 38.220 71.595 ;
        RECT 38.840 70.555 39.010 71.595 ;
        RECT 39.430 70.555 39.600 71.595 ;
        RECT 40.220 70.555 40.390 71.595 ;
        RECT 38.280 69.255 38.780 69.425 ;
        RECT 39.660 69.255 40.160 69.425 ;
        RECT 38.050 68.000 38.220 69.040 ;
        RECT 38.840 68.000 39.010 69.040 ;
        RECT 39.430 68.000 39.600 69.040 ;
        RECT 40.220 68.000 40.390 69.040 ;
        RECT 40.935 67.540 41.645 72.115 ;
        RECT 42.135 67.545 42.845 72.120 ;
        RECT 43.385 70.555 43.555 71.595 ;
        RECT 44.175 70.555 44.345 71.595 ;
        RECT 44.765 70.555 44.935 71.595 ;
        RECT 45.555 70.555 45.725 71.595 ;
        RECT 43.615 69.255 44.115 69.425 ;
        RECT 44.995 69.255 45.495 69.425 ;
        RECT 43.385 68.000 43.555 69.040 ;
        RECT 44.175 68.000 44.345 69.040 ;
        RECT 44.765 68.000 44.935 69.040 ;
        RECT 45.555 68.000 45.725 69.040 ;
        RECT 46.270 67.540 46.980 72.115 ;
        RECT 47.460 67.545 48.170 72.120 ;
        RECT 48.710 70.555 48.880 71.595 ;
        RECT 49.500 70.555 49.670 71.595 ;
        RECT 50.090 70.555 50.260 71.595 ;
        RECT 50.880 70.555 51.050 71.595 ;
        RECT 48.940 69.255 49.440 69.425 ;
        RECT 50.320 69.255 50.820 69.425 ;
        RECT 48.710 68.000 48.880 69.040 ;
        RECT 49.500 68.000 49.670 69.040 ;
        RECT 50.090 68.000 50.260 69.040 ;
        RECT 50.880 68.000 51.050 69.040 ;
        RECT 51.595 67.540 52.305 72.115 ;
        RECT 52.795 67.545 53.505 72.120 ;
        RECT 54.045 70.555 54.215 71.595 ;
        RECT 54.835 70.555 55.005 71.595 ;
        RECT 55.425 70.555 55.595 71.595 ;
        RECT 56.215 70.555 56.385 71.595 ;
        RECT 54.275 69.255 54.775 69.425 ;
        RECT 55.655 69.255 56.155 69.425 ;
        RECT 54.835 68.000 55.005 69.040 ;
        RECT 55.425 68.000 55.595 69.040 ;
        RECT 56.215 68.000 56.385 69.040 ;
        RECT 56.930 67.540 57.640 72.115 ;
        RECT 58.120 67.545 58.830 72.120 ;
        RECT 59.370 70.555 59.540 71.595 ;
        RECT 60.160 70.555 60.330 71.595 ;
        RECT 60.750 70.555 60.920 71.595 ;
        RECT 61.540 70.555 61.710 71.595 ;
        RECT 59.600 69.255 60.100 69.425 ;
        RECT 60.980 69.255 61.480 69.425 ;
        RECT 59.370 68.000 59.540 69.040 ;
        RECT 60.160 68.000 60.330 69.040 ;
        RECT 60.750 68.000 60.920 69.040 ;
        RECT 61.540 68.000 61.710 69.040 ;
        RECT 62.255 67.540 62.965 72.115 ;
        RECT 63.455 67.545 64.165 72.120 ;
        RECT 64.705 70.555 64.875 71.595 ;
        RECT 65.495 70.555 65.665 71.595 ;
        RECT 66.085 70.555 66.255 71.595 ;
        RECT 66.875 70.555 67.045 71.595 ;
        RECT 64.935 69.255 65.435 69.425 ;
        RECT 66.315 69.255 66.815 69.425 ;
        RECT 64.705 68.000 64.875 69.040 ;
        RECT 65.495 68.000 65.665 69.040 ;
        RECT 66.085 68.000 66.255 69.040 ;
        RECT 66.875 68.000 67.045 69.040 ;
        RECT 67.590 67.540 68.300 72.115 ;
        RECT 68.780 67.545 69.490 72.120 ;
        RECT 70.030 70.555 70.200 71.595 ;
        RECT 70.820 70.555 70.990 71.595 ;
        RECT 71.410 70.555 71.580 71.595 ;
        RECT 72.200 70.555 72.370 71.595 ;
        RECT 70.260 69.255 70.760 69.425 ;
        RECT 71.640 69.255 72.140 69.425 ;
        RECT 70.030 68.000 70.200 69.040 ;
        RECT 70.820 68.000 70.990 69.040 ;
        RECT 71.410 68.000 71.580 69.040 ;
        RECT 72.200 68.000 72.370 69.040 ;
        RECT 72.915 67.540 73.625 72.115 ;
        RECT 74.115 67.545 74.825 72.120 ;
        RECT 75.365 70.555 75.535 71.595 ;
        RECT 76.155 70.555 76.325 71.595 ;
        RECT 76.745 70.555 76.915 71.595 ;
        RECT 77.535 70.555 77.705 71.595 ;
        RECT 76.975 69.255 77.475 69.425 ;
        RECT 75.365 68.000 75.535 69.040 ;
        RECT 76.155 68.000 76.325 69.040 ;
        RECT 76.745 68.000 76.915 69.040 ;
        RECT 77.535 68.000 77.705 69.040 ;
        RECT 78.250 67.540 78.960 72.115 ;
        RECT 79.440 67.545 80.150 72.120 ;
        RECT 80.690 70.555 80.860 71.595 ;
        RECT 81.480 70.555 81.650 71.595 ;
        RECT 82.070 70.555 82.240 71.595 ;
        RECT 82.860 70.555 83.030 71.595 ;
        RECT 80.920 69.255 81.420 69.425 ;
        RECT 82.300 69.255 82.800 69.425 ;
        RECT 80.690 68.000 80.860 69.040 ;
        RECT 81.480 68.000 81.650 69.040 ;
        RECT 82.070 68.000 82.240 69.040 ;
        RECT 82.860 68.000 83.030 69.040 ;
        RECT 83.575 67.540 84.285 72.115 ;
        RECT 84.775 67.545 85.485 72.120 ;
        RECT 86.025 70.555 86.195 71.595 ;
        RECT 86.815 70.555 86.985 71.595 ;
        RECT 87.405 70.555 87.575 71.595 ;
        RECT 88.195 70.555 88.365 71.595 ;
        RECT 86.255 69.255 86.755 69.425 ;
        RECT 87.635 69.255 88.135 69.425 ;
        RECT 86.025 68.000 86.195 69.040 ;
        RECT 86.815 68.000 86.985 69.040 ;
        RECT 87.405 68.000 87.575 69.040 ;
        RECT 88.195 68.000 88.365 69.040 ;
        RECT 88.910 67.540 89.620 72.115 ;
        RECT 90.100 67.545 90.810 72.120 ;
        RECT 91.350 70.555 91.520 71.595 ;
        RECT 92.140 70.555 92.310 71.595 ;
        RECT 92.730 70.555 92.900 71.595 ;
        RECT 93.520 70.555 93.690 71.595 ;
        RECT 91.580 69.255 92.080 69.425 ;
        RECT 92.960 69.255 93.460 69.425 ;
        RECT 91.350 68.000 91.520 69.040 ;
        RECT 92.140 68.000 92.310 69.040 ;
        RECT 92.730 68.000 92.900 69.040 ;
        RECT 93.520 68.000 93.690 69.040 ;
        RECT 94.235 67.540 94.945 72.115 ;
        RECT 95.435 67.545 96.145 72.120 ;
        RECT 96.685 70.555 96.855 71.595 ;
        RECT 97.475 70.555 97.645 71.595 ;
        RECT 98.065 70.555 98.235 71.595 ;
        RECT 98.855 70.555 99.025 71.595 ;
        RECT 96.915 69.255 97.415 69.425 ;
        RECT 98.295 69.255 98.795 69.425 ;
        RECT 97.475 68.000 97.645 69.040 ;
        RECT 98.065 68.000 98.235 69.040 ;
        RECT 98.855 68.000 99.025 69.040 ;
        RECT 99.570 67.540 100.280 72.115 ;
        RECT 100.760 67.545 101.470 72.120 ;
        RECT 102.010 70.555 102.180 71.595 ;
        RECT 102.800 70.555 102.970 71.595 ;
        RECT 103.390 70.555 103.560 71.595 ;
        RECT 104.180 70.555 104.350 71.595 ;
        RECT 102.240 69.255 102.740 69.425 ;
        RECT 103.620 69.255 104.120 69.425 ;
        RECT 102.010 68.000 102.180 69.040 ;
        RECT 102.800 68.000 102.970 69.040 ;
        RECT 103.390 68.000 103.560 69.040 ;
        RECT 104.180 68.000 104.350 69.040 ;
        RECT 104.895 67.540 105.605 72.115 ;
        RECT 106.095 67.545 106.805 72.120 ;
        RECT 107.345 70.555 107.515 71.595 ;
        RECT 108.135 70.555 108.305 71.595 ;
        RECT 108.725 70.555 108.895 71.595 ;
        RECT 109.515 70.555 109.685 71.595 ;
        RECT 107.575 69.255 108.075 69.425 ;
        RECT 108.955 69.255 109.455 69.425 ;
        RECT 107.345 68.000 107.515 69.040 ;
        RECT 108.135 68.000 108.305 69.040 ;
        RECT 108.725 68.000 108.895 69.040 ;
        RECT 109.515 68.000 109.685 69.040 ;
        RECT 110.230 67.540 110.940 72.115 ;
        RECT 111.420 67.545 112.130 72.120 ;
        RECT 112.670 70.555 112.840 71.595 ;
        RECT 113.460 70.555 113.630 71.595 ;
        RECT 114.050 70.555 114.220 71.595 ;
        RECT 114.840 70.555 115.010 71.595 ;
        RECT 112.900 69.255 113.400 69.425 ;
        RECT 114.280 69.255 114.780 69.425 ;
        RECT 112.670 68.000 112.840 69.040 ;
        RECT 113.460 68.000 113.630 69.040 ;
        RECT 114.050 68.000 114.220 69.040 ;
        RECT 114.840 68.000 115.010 69.040 ;
        RECT 115.555 67.540 116.265 72.115 ;
        RECT 116.755 67.545 117.465 72.120 ;
        RECT 118.005 70.555 118.175 71.595 ;
        RECT 118.795 70.555 118.965 71.595 ;
        RECT 119.385 70.555 119.555 71.595 ;
        RECT 120.175 70.555 120.345 71.595 ;
        RECT 119.615 69.255 120.115 69.425 ;
        RECT 118.005 68.000 118.175 69.040 ;
        RECT 118.795 68.000 118.965 69.040 ;
        RECT 119.385 68.000 119.555 69.040 ;
        RECT 120.175 68.000 120.345 69.040 ;
        RECT 120.890 67.540 121.600 72.115 ;
        RECT 122.080 67.560 122.790 72.135 ;
        RECT 123.330 70.555 123.500 71.595 ;
        RECT 124.120 70.555 124.290 71.595 ;
        RECT 124.710 70.555 124.880 71.595 ;
        RECT 125.500 70.555 125.670 71.595 ;
        RECT 123.330 68.000 123.500 69.040 ;
        RECT 124.120 68.000 124.290 69.040 ;
        RECT 124.710 68.000 124.880 69.040 ;
        RECT 125.500 68.000 125.670 69.040 ;
        RECT 126.215 67.560 126.925 72.135 ;
        RECT 32.725 66.555 32.895 67.245 ;
        RECT 33.515 66.555 33.685 67.245 ;
        RECT 34.105 66.555 34.275 67.245 ;
        RECT 34.895 66.555 35.065 67.245 ;
        RECT 38.050 66.555 38.220 67.245 ;
        RECT 38.840 66.555 39.010 67.245 ;
        RECT 39.430 66.555 39.600 67.245 ;
        RECT 40.220 66.555 40.390 67.245 ;
        RECT 43.385 66.555 43.555 67.245 ;
        RECT 44.175 66.555 44.345 67.245 ;
        RECT 44.765 66.555 44.935 67.245 ;
        RECT 45.555 66.555 45.725 67.245 ;
        RECT 48.710 66.555 48.880 67.245 ;
        RECT 49.500 66.555 49.670 67.245 ;
        RECT 50.090 66.555 50.260 67.245 ;
        RECT 50.880 66.555 51.050 67.245 ;
        RECT 54.835 66.555 55.005 67.245 ;
        RECT 55.425 66.555 55.595 67.245 ;
        RECT 56.215 66.555 56.385 67.245 ;
        RECT 59.370 66.555 59.540 67.245 ;
        RECT 60.160 66.555 60.330 67.245 ;
        RECT 60.750 66.555 60.920 67.245 ;
        RECT 61.540 66.555 61.710 67.245 ;
        RECT 64.705 66.555 64.875 67.245 ;
        RECT 65.495 66.555 65.665 67.245 ;
        RECT 66.085 66.555 66.255 67.245 ;
        RECT 66.875 66.555 67.045 67.245 ;
        RECT 70.030 66.555 70.200 67.245 ;
        RECT 70.820 66.555 70.990 67.245 ;
        RECT 71.410 66.555 71.580 67.245 ;
        RECT 72.200 66.555 72.370 67.245 ;
        RECT 75.365 66.555 75.535 67.245 ;
        RECT 76.155 66.555 76.325 67.245 ;
        RECT 76.745 66.555 76.915 67.245 ;
        RECT 77.535 66.555 77.705 67.245 ;
        RECT 80.690 66.555 80.860 67.245 ;
        RECT 81.480 66.555 81.650 67.245 ;
        RECT 82.070 66.555 82.240 67.245 ;
        RECT 82.860 66.555 83.030 67.245 ;
        RECT 86.025 66.555 86.195 67.245 ;
        RECT 86.815 66.555 86.985 67.245 ;
        RECT 87.405 66.555 87.575 67.245 ;
        RECT 88.195 66.555 88.365 67.245 ;
        RECT 91.350 66.555 91.520 67.245 ;
        RECT 92.140 66.555 92.310 67.245 ;
        RECT 92.730 66.555 92.900 67.245 ;
        RECT 93.520 66.555 93.690 67.245 ;
        RECT 97.475 66.555 97.645 67.245 ;
        RECT 98.065 66.555 98.235 67.245 ;
        RECT 98.855 66.555 99.025 67.245 ;
        RECT 102.010 66.555 102.180 67.245 ;
        RECT 102.800 66.555 102.970 67.245 ;
        RECT 103.390 66.555 103.560 67.245 ;
        RECT 104.180 66.555 104.350 67.245 ;
        RECT 107.345 66.555 107.515 67.245 ;
        RECT 108.135 66.555 108.305 67.245 ;
        RECT 108.725 66.555 108.895 67.245 ;
        RECT 109.515 66.555 109.685 67.245 ;
        RECT 112.670 66.555 112.840 67.245 ;
        RECT 113.460 66.555 113.630 67.245 ;
        RECT 114.050 66.555 114.220 67.245 ;
        RECT 114.840 66.555 115.010 67.245 ;
        RECT 118.005 66.555 118.175 67.245 ;
        RECT 118.795 66.555 118.965 67.245 ;
        RECT 119.385 66.555 119.555 67.245 ;
        RECT 120.175 66.555 120.345 67.245 ;
        RECT 123.330 66.555 123.500 67.245 ;
        RECT 124.120 66.555 124.290 67.245 ;
        RECT 124.710 66.555 124.880 67.245 ;
        RECT 125.500 66.555 125.670 67.245 ;
        RECT 2.825 64.725 3.155 66.275 ;
        RECT 4.385 64.725 4.715 66.275 ;
        RECT 5.945 64.725 6.275 66.355 ;
        RECT 8.845 65.285 9.175 66.355 ;
        RECT 10.450 65.455 10.780 66.355 ;
        RECT 11.930 65.640 12.180 66.375 ;
        RECT 13.490 65.640 14.075 66.375 ;
        RECT 38.280 66.215 38.780 66.385 ;
        RECT 39.660 66.215 40.160 66.385 ;
        RECT 43.615 66.215 44.115 66.385 ;
        RECT 44.995 66.215 45.495 66.385 ;
        RECT 48.940 66.215 49.440 66.385 ;
        RECT 50.320 66.215 50.820 66.385 ;
        RECT 54.275 66.215 54.775 66.385 ;
        RECT 55.655 66.215 56.155 66.385 ;
        RECT 59.600 66.215 60.100 66.385 ;
        RECT 60.980 66.215 61.480 66.385 ;
        RECT 64.935 66.215 65.435 66.385 ;
        RECT 66.315 66.215 66.815 66.385 ;
        RECT 70.260 66.215 70.760 66.385 ;
        RECT 71.640 66.215 72.140 66.385 ;
        RECT 76.975 66.215 77.475 66.385 ;
        RECT 80.920 66.215 81.420 66.385 ;
        RECT 82.300 66.215 82.800 66.385 ;
        RECT 86.255 66.215 86.755 66.385 ;
        RECT 87.635 66.215 88.135 66.385 ;
        RECT 91.580 66.215 92.080 66.385 ;
        RECT 92.960 66.215 93.460 66.385 ;
        RECT 96.915 66.215 97.415 66.385 ;
        RECT 98.295 66.215 98.795 66.385 ;
        RECT 102.240 66.215 102.740 66.385 ;
        RECT 103.620 66.215 104.120 66.385 ;
        RECT 107.575 66.215 108.075 66.385 ;
        RECT 108.955 66.215 109.455 66.385 ;
        RECT 112.900 66.215 113.400 66.385 ;
        RECT 114.280 66.215 114.780 66.385 ;
        RECT 119.615 66.215 120.115 66.385 ;
        RECT 11.930 65.470 14.075 65.640 ;
        RECT 15.925 65.645 16.135 66.140 ;
        RECT 17.485 65.645 17.695 66.140 ;
        RECT 19.045 65.645 19.255 66.140 ;
        RECT 20.645 65.645 21.295 66.140 ;
        RECT 38.280 65.675 38.780 65.845 ;
        RECT 39.660 65.675 40.160 65.845 ;
        RECT 43.615 65.675 44.115 65.845 ;
        RECT 44.995 65.675 45.495 65.845 ;
        RECT 48.940 65.675 49.440 65.845 ;
        RECT 50.320 65.675 50.820 65.845 ;
        RECT 54.275 65.675 54.775 65.845 ;
        RECT 55.655 65.675 56.155 65.845 ;
        RECT 59.600 65.675 60.100 65.845 ;
        RECT 60.980 65.675 61.480 65.845 ;
        RECT 64.935 65.675 65.435 65.845 ;
        RECT 66.315 65.675 66.815 65.845 ;
        RECT 70.260 65.675 70.760 65.845 ;
        RECT 71.640 65.675 72.140 65.845 ;
        RECT 75.595 65.675 76.095 65.845 ;
        RECT 76.975 65.675 77.475 65.845 ;
        RECT 80.920 65.675 81.420 65.845 ;
        RECT 82.300 65.675 82.800 65.845 ;
        RECT 86.255 65.675 86.755 65.845 ;
        RECT 87.635 65.675 88.135 65.845 ;
        RECT 91.580 65.675 92.080 65.845 ;
        RECT 92.960 65.675 93.460 65.845 ;
        RECT 96.915 65.675 97.415 65.845 ;
        RECT 98.295 65.675 98.795 65.845 ;
        RECT 102.240 65.675 102.740 65.845 ;
        RECT 103.620 65.675 104.120 65.845 ;
        RECT 107.575 65.675 108.075 65.845 ;
        RECT 108.955 65.675 109.455 65.845 ;
        RECT 112.900 65.675 113.400 65.845 ;
        RECT 114.280 65.675 114.780 65.845 ;
        RECT 118.235 65.675 118.735 65.845 ;
        RECT 119.615 65.675 120.115 65.845 ;
        RECT 15.925 65.470 21.840 65.645 ;
        RECT 7.990 64.725 8.320 65.285 ;
        RECT 2.825 64.395 8.320 64.725 ;
        RECT 3.215 61.785 3.505 64.225 ;
        RECT 6.515 62.195 6.845 64.395 ;
        RECT 7.990 63.935 8.320 64.395 ;
        RECT 8.845 64.955 10.370 65.285 ;
        RECT 7.015 63.200 7.825 63.530 ;
        RECT 7.495 62.535 7.825 63.200 ;
        RECT 8.845 63.135 9.175 64.955 ;
        RECT 10.540 64.785 10.780 65.455 ;
        RECT 13.905 65.320 14.075 65.470 ;
        RECT 13.905 65.290 14.605 65.320 ;
        RECT 11.015 65.120 13.725 65.290 ;
        RECT 13.905 65.055 21.490 65.290 ;
        RECT 13.905 64.940 15.710 65.055 ;
        RECT 10.450 63.135 10.780 64.785 ;
        RECT 11.930 64.770 15.710 64.940 ;
        RECT 21.670 64.840 21.840 65.470 ;
        RECT 16.045 64.835 21.840 64.840 ;
        RECT 11.930 63.115 12.260 64.770 ;
        RECT 13.570 63.115 13.820 64.770 ;
        RECT 16.005 64.665 21.840 64.835 ;
        RECT 32.725 64.815 32.895 65.505 ;
        RECT 33.515 64.815 33.685 65.505 ;
        RECT 34.105 64.815 34.275 65.505 ;
        RECT 34.895 64.815 35.065 65.505 ;
        RECT 38.050 64.815 38.220 65.505 ;
        RECT 38.840 64.815 39.010 65.505 ;
        RECT 39.430 64.815 39.600 65.505 ;
        RECT 40.220 64.815 40.390 65.505 ;
        RECT 43.385 64.815 43.555 65.505 ;
        RECT 44.175 64.815 44.345 65.505 ;
        RECT 44.765 64.815 44.935 65.505 ;
        RECT 45.555 64.815 45.725 65.505 ;
        RECT 48.710 64.815 48.880 65.505 ;
        RECT 49.500 64.815 49.670 65.505 ;
        RECT 50.090 64.815 50.260 65.505 ;
        RECT 50.880 64.815 51.050 65.505 ;
        RECT 54.045 64.815 54.215 65.505 ;
        RECT 54.835 64.815 55.005 65.505 ;
        RECT 55.425 64.815 55.595 65.505 ;
        RECT 56.215 64.815 56.385 65.505 ;
        RECT 59.370 64.815 59.540 65.505 ;
        RECT 60.160 64.815 60.330 65.505 ;
        RECT 60.750 64.815 60.920 65.505 ;
        RECT 61.540 64.815 61.710 65.505 ;
        RECT 64.705 64.815 64.875 65.505 ;
        RECT 65.495 64.815 65.665 65.505 ;
        RECT 66.085 64.815 66.255 65.505 ;
        RECT 66.875 64.815 67.045 65.505 ;
        RECT 70.030 64.815 70.200 65.505 ;
        RECT 70.820 64.815 70.990 65.505 ;
        RECT 71.410 64.815 71.580 65.505 ;
        RECT 72.200 64.815 72.370 65.505 ;
        RECT 75.365 64.815 75.535 65.505 ;
        RECT 76.155 64.815 76.325 65.505 ;
        RECT 76.745 64.815 76.915 65.505 ;
        RECT 77.535 64.815 77.705 65.505 ;
        RECT 80.690 64.815 80.860 65.505 ;
        RECT 81.480 64.815 81.650 65.505 ;
        RECT 82.070 64.815 82.240 65.505 ;
        RECT 82.860 64.815 83.030 65.505 ;
        RECT 86.025 64.815 86.195 65.505 ;
        RECT 86.815 64.815 86.985 65.505 ;
        RECT 87.405 64.815 87.575 65.505 ;
        RECT 88.195 64.815 88.365 65.505 ;
        RECT 91.350 64.815 91.520 65.505 ;
        RECT 92.140 64.815 92.310 65.505 ;
        RECT 92.730 64.815 92.900 65.505 ;
        RECT 93.520 64.815 93.690 65.505 ;
        RECT 96.685 64.815 96.855 65.505 ;
        RECT 97.475 64.815 97.645 65.505 ;
        RECT 98.065 64.815 98.235 65.505 ;
        RECT 98.855 64.815 99.025 65.505 ;
        RECT 102.010 64.815 102.180 65.505 ;
        RECT 102.800 64.815 102.970 65.505 ;
        RECT 103.390 64.815 103.560 65.505 ;
        RECT 104.180 64.815 104.350 65.505 ;
        RECT 107.345 64.815 107.515 65.505 ;
        RECT 108.135 64.815 108.305 65.505 ;
        RECT 108.725 64.815 108.895 65.505 ;
        RECT 109.515 64.815 109.685 65.505 ;
        RECT 112.670 64.815 112.840 65.505 ;
        RECT 113.460 64.815 113.630 65.505 ;
        RECT 114.050 64.815 114.220 65.505 ;
        RECT 114.840 64.815 115.010 65.505 ;
        RECT 118.005 64.815 118.175 65.505 ;
        RECT 118.795 64.815 118.965 65.505 ;
        RECT 119.385 64.815 119.555 65.505 ;
        RECT 120.175 64.815 120.345 65.505 ;
        RECT 123.330 64.815 123.500 65.505 ;
        RECT 124.120 64.815 124.290 65.505 ;
        RECT 124.710 64.815 124.880 65.505 ;
        RECT 125.500 64.815 125.670 65.505 ;
        RECT 16.005 63.425 16.335 64.665 ;
        RECT 17.565 63.425 17.895 64.665 ;
        RECT 19.125 63.425 19.455 64.665 ;
        RECT 20.685 63.425 21.015 64.665 ;
        RECT 6.515 61.865 7.325 62.195 ;
        RECT 3.215 61.495 3.595 61.785 ;
        RECT 3.305 60.725 3.595 61.495 ;
        RECT 4.205 61.205 4.515 61.635 ;
        RECT 6.995 61.525 7.325 61.865 ;
        RECT 7.495 62.125 8.165 62.535 ;
        RECT 7.495 61.205 7.825 62.125 ;
        RECT 4.205 60.895 6.120 61.205 ;
        RECT 4.810 60.875 6.120 60.895 ;
        RECT 6.290 60.875 9.740 61.205 ;
        RECT 3.305 60.475 4.640 60.725 ;
        RECT 3.305 59.465 3.595 60.475 ;
        RECT 4.810 60.305 5.140 60.875 ;
        RECT 4.205 59.975 5.140 60.305 ;
        RECT 4.205 59.465 4.515 59.975 ;
        RECT 6.290 59.325 6.620 60.875 ;
        RECT 7.850 59.325 8.180 60.875 ;
        RECT 9.410 59.245 9.740 60.875 ;
        RECT 11.015 60.280 11.960 60.610 ;
        RECT 12.130 60.510 12.380 62.485 ;
        RECT 14.565 60.935 14.895 62.175 ;
        RECT 16.125 60.935 16.455 62.175 ;
        RECT 17.685 60.935 18.015 62.175 ;
        RECT 19.245 60.935 19.575 62.175 ;
        RECT 14.565 60.765 20.400 60.935 ;
        RECT 16.175 60.750 20.400 60.765 ;
        RECT 14.645 60.545 15.945 60.575 ;
        RECT 12.130 60.340 12.685 60.510 ;
        RECT 12.455 60.100 12.685 60.340 ;
        RECT 13.600 60.310 20.050 60.545 ;
        RECT 12.090 59.270 12.685 60.100 ;
        RECT 14.485 60.125 19.515 60.130 ;
        RECT 20.230 60.125 20.400 60.750 ;
        RECT 14.485 59.960 20.400 60.125 ;
        RECT 31.475 60.025 32.185 64.600 ;
        RECT 32.725 63.020 32.895 64.060 ;
        RECT 33.515 63.020 33.685 64.060 ;
        RECT 34.105 63.020 34.275 64.060 ;
        RECT 34.895 63.020 35.065 64.060 ;
        RECT 32.725 60.465 32.895 61.505 ;
        RECT 33.515 60.465 33.685 61.505 ;
        RECT 34.105 60.465 34.275 61.505 ;
        RECT 34.895 60.465 35.065 61.505 ;
        RECT 35.610 60.025 36.320 64.600 ;
        RECT 36.800 60.010 37.510 64.585 ;
        RECT 38.050 63.020 38.220 64.060 ;
        RECT 38.840 63.020 39.010 64.060 ;
        RECT 39.430 63.020 39.600 64.060 ;
        RECT 40.220 63.020 40.390 64.060 ;
        RECT 38.280 62.635 38.780 62.805 ;
        RECT 39.660 62.635 40.160 62.805 ;
        RECT 38.280 61.720 38.780 61.890 ;
        RECT 39.660 61.720 40.160 61.890 ;
        RECT 38.050 60.465 38.220 61.505 ;
        RECT 38.840 60.465 39.010 61.505 ;
        RECT 39.430 60.465 39.600 61.505 ;
        RECT 40.220 60.465 40.390 61.505 ;
        RECT 40.935 60.005 41.645 64.580 ;
        RECT 42.135 60.010 42.845 64.585 ;
        RECT 43.385 63.020 43.555 64.060 ;
        RECT 44.175 63.020 44.345 64.060 ;
        RECT 44.765 63.020 44.935 64.060 ;
        RECT 45.555 63.020 45.725 64.060 ;
        RECT 43.615 62.635 44.115 62.805 ;
        RECT 44.995 62.635 45.495 62.805 ;
        RECT 43.615 61.720 44.115 61.890 ;
        RECT 44.995 61.720 45.495 61.890 ;
        RECT 43.385 60.465 43.555 61.505 ;
        RECT 44.175 60.465 44.345 61.505 ;
        RECT 44.765 60.465 44.935 61.505 ;
        RECT 45.555 60.465 45.725 61.505 ;
        RECT 46.270 60.005 46.980 64.580 ;
        RECT 47.460 60.010 48.170 64.585 ;
        RECT 48.710 63.020 48.880 64.060 ;
        RECT 49.500 63.020 49.670 64.060 ;
        RECT 50.090 63.020 50.260 64.060 ;
        RECT 50.880 63.020 51.050 64.060 ;
        RECT 48.940 62.635 49.440 62.805 ;
        RECT 50.320 62.635 50.820 62.805 ;
        RECT 48.940 61.720 49.440 61.890 ;
        RECT 50.320 61.720 50.820 61.890 ;
        RECT 48.710 60.465 48.880 61.505 ;
        RECT 49.500 60.465 49.670 61.505 ;
        RECT 50.090 60.465 50.260 61.505 ;
        RECT 50.880 60.465 51.050 61.505 ;
        RECT 51.595 60.005 52.305 64.580 ;
        RECT 52.795 60.010 53.505 64.585 ;
        RECT 54.045 63.020 54.215 64.060 ;
        RECT 54.835 63.020 55.005 64.060 ;
        RECT 55.425 63.020 55.595 64.060 ;
        RECT 56.215 63.020 56.385 64.060 ;
        RECT 54.275 62.635 54.775 62.805 ;
        RECT 55.655 62.635 56.155 62.805 ;
        RECT 54.275 61.720 54.775 61.890 ;
        RECT 55.655 61.720 56.155 61.890 ;
        RECT 54.045 60.465 54.215 61.505 ;
        RECT 54.835 60.465 55.005 61.505 ;
        RECT 55.425 60.465 55.595 61.505 ;
        RECT 56.215 60.465 56.385 61.505 ;
        RECT 56.930 60.005 57.640 64.580 ;
        RECT 58.120 60.010 58.830 64.585 ;
        RECT 59.370 63.020 59.540 64.060 ;
        RECT 60.160 63.020 60.330 64.060 ;
        RECT 60.750 63.020 60.920 64.060 ;
        RECT 61.540 63.020 61.710 64.060 ;
        RECT 59.600 62.635 60.100 62.805 ;
        RECT 60.980 62.635 61.480 62.805 ;
        RECT 59.600 61.720 60.100 61.890 ;
        RECT 60.980 61.720 61.480 61.890 ;
        RECT 59.370 60.465 59.540 61.505 ;
        RECT 60.160 60.465 60.330 61.505 ;
        RECT 60.750 60.465 60.920 61.505 ;
        RECT 61.540 60.465 61.710 61.505 ;
        RECT 62.255 60.005 62.965 64.580 ;
        RECT 63.455 60.010 64.165 64.585 ;
        RECT 64.705 63.020 64.875 64.060 ;
        RECT 65.495 63.020 65.665 64.060 ;
        RECT 66.085 63.020 66.255 64.060 ;
        RECT 66.875 63.020 67.045 64.060 ;
        RECT 64.935 62.635 65.435 62.805 ;
        RECT 66.315 62.635 66.815 62.805 ;
        RECT 64.935 61.720 65.435 61.890 ;
        RECT 66.315 61.720 66.815 61.890 ;
        RECT 64.705 60.465 64.875 61.505 ;
        RECT 65.495 60.465 65.665 61.505 ;
        RECT 66.085 60.465 66.255 61.505 ;
        RECT 66.875 60.465 67.045 61.505 ;
        RECT 67.590 60.005 68.300 64.580 ;
        RECT 68.780 60.010 69.490 64.585 ;
        RECT 70.030 63.020 70.200 64.060 ;
        RECT 70.820 63.020 70.990 64.060 ;
        RECT 71.410 63.020 71.580 64.060 ;
        RECT 72.200 63.020 72.370 64.060 ;
        RECT 70.260 62.635 70.760 62.805 ;
        RECT 71.640 62.635 72.140 62.805 ;
        RECT 70.260 61.720 70.760 61.890 ;
        RECT 71.640 61.720 72.140 61.890 ;
        RECT 70.030 60.465 70.200 61.505 ;
        RECT 70.820 60.465 70.990 61.505 ;
        RECT 71.410 60.465 71.580 61.505 ;
        RECT 72.200 60.465 72.370 61.505 ;
        RECT 72.915 60.005 73.625 64.580 ;
        RECT 74.115 60.010 74.825 64.585 ;
        RECT 75.365 63.020 75.535 64.060 ;
        RECT 76.155 63.020 76.325 64.060 ;
        RECT 76.745 63.020 76.915 64.060 ;
        RECT 77.535 63.020 77.705 64.060 ;
        RECT 75.595 62.635 76.095 62.805 ;
        RECT 76.975 62.635 77.475 62.805 ;
        RECT 75.595 61.720 76.095 61.890 ;
        RECT 76.975 61.720 77.475 61.890 ;
        RECT 75.365 60.465 75.535 61.505 ;
        RECT 76.155 60.465 76.325 61.505 ;
        RECT 76.745 60.465 76.915 61.505 ;
        RECT 77.535 60.465 77.705 61.505 ;
        RECT 78.250 60.005 78.960 64.580 ;
        RECT 79.440 60.010 80.150 64.585 ;
        RECT 80.690 63.020 80.860 64.060 ;
        RECT 81.480 63.020 81.650 64.060 ;
        RECT 82.070 63.020 82.240 64.060 ;
        RECT 82.860 63.020 83.030 64.060 ;
        RECT 80.920 62.635 81.420 62.805 ;
        RECT 82.300 62.635 82.800 62.805 ;
        RECT 80.920 61.720 81.420 61.890 ;
        RECT 82.300 61.720 82.800 61.890 ;
        RECT 80.690 60.465 80.860 61.505 ;
        RECT 81.480 60.465 81.650 61.505 ;
        RECT 82.070 60.465 82.240 61.505 ;
        RECT 82.860 60.465 83.030 61.505 ;
        RECT 83.575 60.005 84.285 64.580 ;
        RECT 84.775 60.010 85.485 64.585 ;
        RECT 86.025 63.020 86.195 64.060 ;
        RECT 86.815 63.020 86.985 64.060 ;
        RECT 87.405 63.020 87.575 64.060 ;
        RECT 88.195 63.020 88.365 64.060 ;
        RECT 86.255 62.635 86.755 62.805 ;
        RECT 87.635 62.635 88.135 62.805 ;
        RECT 86.255 61.720 86.755 61.890 ;
        RECT 87.635 61.720 88.135 61.890 ;
        RECT 86.025 60.465 86.195 61.505 ;
        RECT 86.815 60.465 86.985 61.505 ;
        RECT 87.405 60.465 87.575 61.505 ;
        RECT 88.195 60.465 88.365 61.505 ;
        RECT 88.910 60.005 89.620 64.580 ;
        RECT 90.100 60.010 90.810 64.585 ;
        RECT 91.350 63.020 91.520 64.060 ;
        RECT 92.140 63.020 92.310 64.060 ;
        RECT 92.730 63.020 92.900 64.060 ;
        RECT 93.520 63.020 93.690 64.060 ;
        RECT 91.580 62.635 92.080 62.805 ;
        RECT 92.960 62.635 93.460 62.805 ;
        RECT 91.580 61.720 92.080 61.890 ;
        RECT 92.960 61.720 93.460 61.890 ;
        RECT 91.350 60.465 91.520 61.505 ;
        RECT 92.140 60.465 92.310 61.505 ;
        RECT 92.730 60.465 92.900 61.505 ;
        RECT 93.520 60.465 93.690 61.505 ;
        RECT 94.235 60.005 94.945 64.580 ;
        RECT 95.435 60.010 96.145 64.585 ;
        RECT 96.685 63.020 96.855 64.060 ;
        RECT 97.475 63.020 97.645 64.060 ;
        RECT 98.065 63.020 98.235 64.060 ;
        RECT 98.855 63.020 99.025 64.060 ;
        RECT 96.915 62.635 97.415 62.805 ;
        RECT 98.295 62.635 98.795 62.805 ;
        RECT 96.915 61.720 97.415 61.890 ;
        RECT 98.295 61.720 98.795 61.890 ;
        RECT 96.685 60.465 96.855 61.505 ;
        RECT 97.475 60.465 97.645 61.505 ;
        RECT 98.065 60.465 98.235 61.505 ;
        RECT 98.855 60.465 99.025 61.505 ;
        RECT 99.570 60.005 100.280 64.580 ;
        RECT 100.760 60.010 101.470 64.585 ;
        RECT 102.010 63.020 102.180 64.060 ;
        RECT 102.800 63.020 102.970 64.060 ;
        RECT 103.390 63.020 103.560 64.060 ;
        RECT 104.180 63.020 104.350 64.060 ;
        RECT 102.240 62.635 102.740 62.805 ;
        RECT 103.620 62.635 104.120 62.805 ;
        RECT 102.240 61.720 102.740 61.890 ;
        RECT 103.620 61.720 104.120 61.890 ;
        RECT 102.010 60.465 102.180 61.505 ;
        RECT 102.800 60.465 102.970 61.505 ;
        RECT 103.390 60.465 103.560 61.505 ;
        RECT 104.180 60.465 104.350 61.505 ;
        RECT 104.895 60.005 105.605 64.580 ;
        RECT 106.095 60.010 106.805 64.585 ;
        RECT 107.345 63.020 107.515 64.060 ;
        RECT 108.135 63.020 108.305 64.060 ;
        RECT 108.725 63.020 108.895 64.060 ;
        RECT 109.515 63.020 109.685 64.060 ;
        RECT 107.575 62.635 108.075 62.805 ;
        RECT 108.955 62.635 109.455 62.805 ;
        RECT 107.575 61.720 108.075 61.890 ;
        RECT 108.955 61.720 109.455 61.890 ;
        RECT 107.345 60.465 107.515 61.505 ;
        RECT 108.135 60.465 108.305 61.505 ;
        RECT 108.725 60.465 108.895 61.505 ;
        RECT 109.515 60.465 109.685 61.505 ;
        RECT 110.230 60.005 110.940 64.580 ;
        RECT 111.420 60.010 112.130 64.585 ;
        RECT 112.670 63.020 112.840 64.060 ;
        RECT 113.460 63.020 113.630 64.060 ;
        RECT 114.050 63.020 114.220 64.060 ;
        RECT 114.840 63.020 115.010 64.060 ;
        RECT 112.900 62.635 113.400 62.805 ;
        RECT 114.280 62.635 114.780 62.805 ;
        RECT 112.900 61.720 113.400 61.890 ;
        RECT 114.280 61.720 114.780 61.890 ;
        RECT 112.670 60.465 112.840 61.505 ;
        RECT 113.460 60.465 113.630 61.505 ;
        RECT 114.050 60.465 114.220 61.505 ;
        RECT 114.840 60.465 115.010 61.505 ;
        RECT 115.555 60.005 116.265 64.580 ;
        RECT 116.755 60.010 117.465 64.585 ;
        RECT 118.005 63.020 118.175 64.060 ;
        RECT 118.795 63.020 118.965 64.060 ;
        RECT 119.385 63.020 119.555 64.060 ;
        RECT 120.175 63.020 120.345 64.060 ;
        RECT 118.235 62.635 118.735 62.805 ;
        RECT 119.615 62.635 120.115 62.805 ;
        RECT 118.235 61.720 118.735 61.890 ;
        RECT 119.615 61.720 120.115 61.890 ;
        RECT 118.005 60.465 118.175 61.505 ;
        RECT 118.795 60.465 118.965 61.505 ;
        RECT 119.385 60.465 119.555 61.505 ;
        RECT 120.175 60.465 120.345 61.505 ;
        RECT 120.890 60.005 121.600 64.580 ;
        RECT 122.080 60.025 122.790 64.600 ;
        RECT 123.330 63.020 123.500 64.060 ;
        RECT 124.120 63.020 124.290 64.060 ;
        RECT 124.710 63.020 124.880 64.060 ;
        RECT 125.500 63.020 125.670 64.060 ;
        RECT 123.330 60.465 123.500 61.505 ;
        RECT 124.120 60.465 124.290 61.505 ;
        RECT 124.710 60.465 124.880 61.505 ;
        RECT 125.500 60.465 125.670 61.505 ;
        RECT 126.215 60.025 126.925 64.600 ;
        RECT 14.485 59.460 14.695 59.960 ;
        RECT 16.045 59.955 20.400 59.960 ;
        RECT 16.045 59.945 20.260 59.955 ;
        RECT 16.045 59.460 16.255 59.945 ;
        RECT 17.605 59.460 17.815 59.945 ;
        RECT 19.205 59.460 19.855 59.945 ;
        RECT 32.725 59.020 32.895 59.710 ;
        RECT 33.515 59.020 33.685 59.710 ;
        RECT 34.105 59.020 34.275 59.710 ;
        RECT 34.895 59.020 35.065 59.710 ;
        RECT 38.050 59.020 38.220 59.710 ;
        RECT 38.840 59.020 39.010 59.710 ;
        RECT 39.430 59.020 39.600 59.710 ;
        RECT 40.220 59.020 40.390 59.710 ;
        RECT 43.385 59.020 43.555 59.710 ;
        RECT 44.175 59.020 44.345 59.710 ;
        RECT 44.765 59.020 44.935 59.710 ;
        RECT 45.555 59.020 45.725 59.710 ;
        RECT 48.710 59.020 48.880 59.710 ;
        RECT 49.500 59.020 49.670 59.710 ;
        RECT 50.090 59.020 50.260 59.710 ;
        RECT 50.880 59.020 51.050 59.710 ;
        RECT 54.045 59.020 54.215 59.710 ;
        RECT 54.835 59.020 55.005 59.710 ;
        RECT 55.425 59.020 55.595 59.710 ;
        RECT 56.215 59.020 56.385 59.710 ;
        RECT 59.370 59.020 59.540 59.710 ;
        RECT 60.160 59.020 60.330 59.710 ;
        RECT 60.750 59.020 60.920 59.710 ;
        RECT 61.540 59.020 61.710 59.710 ;
        RECT 64.705 59.020 64.875 59.710 ;
        RECT 65.495 59.020 65.665 59.710 ;
        RECT 66.085 59.020 66.255 59.710 ;
        RECT 66.875 59.020 67.045 59.710 ;
        RECT 70.030 59.020 70.200 59.710 ;
        RECT 70.820 59.020 70.990 59.710 ;
        RECT 71.410 59.020 71.580 59.710 ;
        RECT 72.200 59.020 72.370 59.710 ;
        RECT 75.365 59.020 75.535 59.710 ;
        RECT 76.155 59.020 76.325 59.710 ;
        RECT 76.745 59.020 76.915 59.710 ;
        RECT 77.535 59.020 77.705 59.710 ;
        RECT 80.690 59.020 80.860 59.710 ;
        RECT 81.480 59.020 81.650 59.710 ;
        RECT 82.070 59.020 82.240 59.710 ;
        RECT 82.860 59.020 83.030 59.710 ;
        RECT 86.025 59.020 86.195 59.710 ;
        RECT 86.815 59.020 86.985 59.710 ;
        RECT 87.405 59.020 87.575 59.710 ;
        RECT 88.195 59.020 88.365 59.710 ;
        RECT 91.350 59.020 91.520 59.710 ;
        RECT 92.140 59.020 92.310 59.710 ;
        RECT 92.730 59.020 92.900 59.710 ;
        RECT 93.520 59.020 93.690 59.710 ;
        RECT 96.685 59.020 96.855 59.710 ;
        RECT 97.475 59.020 97.645 59.710 ;
        RECT 98.065 59.020 98.235 59.710 ;
        RECT 98.855 59.020 99.025 59.710 ;
        RECT 102.010 59.020 102.180 59.710 ;
        RECT 102.800 59.020 102.970 59.710 ;
        RECT 103.390 59.020 103.560 59.710 ;
        RECT 104.180 59.020 104.350 59.710 ;
        RECT 107.345 59.020 107.515 59.710 ;
        RECT 108.135 59.020 108.305 59.710 ;
        RECT 108.725 59.020 108.895 59.710 ;
        RECT 109.515 59.020 109.685 59.710 ;
        RECT 112.670 59.020 112.840 59.710 ;
        RECT 113.460 59.020 113.630 59.710 ;
        RECT 114.050 59.020 114.220 59.710 ;
        RECT 114.840 59.020 115.010 59.710 ;
        RECT 118.005 59.020 118.175 59.710 ;
        RECT 118.795 59.020 118.965 59.710 ;
        RECT 119.385 59.020 119.555 59.710 ;
        RECT 120.175 59.020 120.345 59.710 ;
        RECT 123.330 59.020 123.500 59.710 ;
        RECT 124.120 59.020 124.290 59.710 ;
        RECT 124.710 59.020 124.880 59.710 ;
        RECT 125.500 59.020 125.670 59.710 ;
        RECT 38.280 58.680 38.780 58.850 ;
        RECT 39.660 58.680 40.160 58.850 ;
        RECT 43.615 58.680 44.115 58.850 ;
        RECT 44.995 58.680 45.495 58.850 ;
        RECT 48.940 58.680 49.440 58.850 ;
        RECT 50.320 58.680 50.820 58.850 ;
        RECT 54.275 58.680 54.775 58.850 ;
        RECT 55.655 58.680 56.155 58.850 ;
        RECT 59.600 58.680 60.100 58.850 ;
        RECT 60.980 58.680 61.480 58.850 ;
        RECT 64.935 58.680 65.435 58.850 ;
        RECT 66.315 58.680 66.815 58.850 ;
        RECT 70.260 58.680 70.760 58.850 ;
        RECT 71.640 58.680 72.140 58.850 ;
        RECT 75.595 58.680 76.095 58.850 ;
        RECT 76.975 58.680 77.475 58.850 ;
        RECT 80.920 58.680 81.420 58.850 ;
        RECT 82.300 58.680 82.800 58.850 ;
        RECT 86.255 58.680 86.755 58.850 ;
        RECT 87.635 58.680 88.135 58.850 ;
        RECT 91.580 58.680 92.080 58.850 ;
        RECT 92.960 58.680 93.460 58.850 ;
        RECT 96.915 58.680 97.415 58.850 ;
        RECT 98.295 58.680 98.795 58.850 ;
        RECT 102.240 58.680 102.740 58.850 ;
        RECT 103.620 58.680 104.120 58.850 ;
        RECT 107.575 58.680 108.075 58.850 ;
        RECT 108.955 58.680 109.455 58.850 ;
        RECT 112.900 58.680 113.400 58.850 ;
        RECT 114.280 58.680 114.780 58.850 ;
        RECT 118.235 58.680 118.735 58.850 ;
        RECT 119.615 58.680 120.115 58.850 ;
        RECT 2.825 56.585 3.155 58.135 ;
        RECT 4.385 56.585 4.715 58.135 ;
        RECT 5.945 56.585 6.275 58.215 ;
        RECT 8.845 57.145 9.175 58.215 ;
        RECT 10.450 57.315 10.780 58.215 ;
        RECT 11.930 57.500 12.180 58.235 ;
        RECT 13.490 57.500 14.075 58.235 ;
        RECT 38.280 58.140 38.780 58.310 ;
        RECT 39.660 58.140 40.160 58.310 ;
        RECT 43.615 58.140 44.115 58.310 ;
        RECT 44.995 58.140 45.495 58.310 ;
        RECT 48.940 58.140 49.440 58.310 ;
        RECT 50.320 58.140 50.820 58.310 ;
        RECT 54.275 58.140 54.775 58.310 ;
        RECT 55.655 58.140 56.155 58.310 ;
        RECT 59.600 58.140 60.100 58.310 ;
        RECT 60.980 58.140 61.480 58.310 ;
        RECT 64.935 58.140 65.435 58.310 ;
        RECT 66.315 58.140 66.815 58.310 ;
        RECT 70.260 58.140 70.760 58.310 ;
        RECT 71.640 58.140 72.140 58.310 ;
        RECT 75.595 58.140 76.095 58.310 ;
        RECT 76.975 58.140 77.475 58.310 ;
        RECT 80.920 58.140 81.420 58.310 ;
        RECT 82.300 58.140 82.800 58.310 ;
        RECT 86.255 58.140 86.755 58.310 ;
        RECT 87.635 58.140 88.135 58.310 ;
        RECT 91.580 58.140 92.080 58.310 ;
        RECT 92.960 58.140 93.460 58.310 ;
        RECT 96.915 58.140 97.415 58.310 ;
        RECT 98.295 58.140 98.795 58.310 ;
        RECT 102.240 58.140 102.740 58.310 ;
        RECT 103.620 58.140 104.120 58.310 ;
        RECT 107.575 58.140 108.075 58.310 ;
        RECT 108.955 58.140 109.455 58.310 ;
        RECT 112.900 58.140 113.400 58.310 ;
        RECT 114.280 58.140 114.780 58.310 ;
        RECT 118.235 58.140 118.735 58.310 ;
        RECT 119.615 58.140 120.115 58.310 ;
        RECT 11.930 57.330 14.075 57.500 ;
        RECT 15.925 57.505 16.135 58.000 ;
        RECT 17.485 57.505 17.695 58.000 ;
        RECT 19.045 57.505 19.255 58.000 ;
        RECT 20.645 57.505 21.295 58.000 ;
        RECT 15.925 57.330 21.840 57.505 ;
        RECT 7.990 56.585 8.320 57.145 ;
        RECT 2.825 56.255 8.320 56.585 ;
        RECT 3.215 53.645 3.505 56.085 ;
        RECT 6.515 54.055 6.845 56.255 ;
        RECT 7.990 55.795 8.320 56.255 ;
        RECT 8.845 56.815 10.370 57.145 ;
        RECT 7.015 55.060 7.825 55.390 ;
        RECT 7.495 54.395 7.825 55.060 ;
        RECT 8.845 54.995 9.175 56.815 ;
        RECT 10.540 56.645 10.780 57.315 ;
        RECT 13.905 57.180 14.075 57.330 ;
        RECT 13.905 57.150 14.605 57.180 ;
        RECT 11.015 56.980 13.725 57.150 ;
        RECT 13.905 56.915 21.490 57.150 ;
        RECT 13.905 56.800 15.710 56.915 ;
        RECT 10.450 54.995 10.780 56.645 ;
        RECT 11.930 56.630 15.710 56.800 ;
        RECT 21.670 56.700 21.840 57.330 ;
        RECT 32.725 57.280 32.895 57.970 ;
        RECT 33.515 57.280 33.685 57.970 ;
        RECT 34.105 57.280 34.275 57.970 ;
        RECT 34.895 57.280 35.065 57.970 ;
        RECT 38.050 57.280 38.220 57.970 ;
        RECT 38.840 57.280 39.010 57.970 ;
        RECT 39.430 57.280 39.600 57.970 ;
        RECT 40.220 57.280 40.390 57.970 ;
        RECT 43.385 57.280 43.555 57.970 ;
        RECT 44.175 57.280 44.345 57.970 ;
        RECT 44.765 57.280 44.935 57.970 ;
        RECT 45.555 57.280 45.725 57.970 ;
        RECT 48.710 57.280 48.880 57.970 ;
        RECT 49.500 57.280 49.670 57.970 ;
        RECT 50.090 57.280 50.260 57.970 ;
        RECT 50.880 57.280 51.050 57.970 ;
        RECT 54.045 57.280 54.215 57.970 ;
        RECT 54.835 57.280 55.005 57.970 ;
        RECT 55.425 57.280 55.595 57.970 ;
        RECT 56.215 57.280 56.385 57.970 ;
        RECT 59.370 57.280 59.540 57.970 ;
        RECT 60.160 57.280 60.330 57.970 ;
        RECT 60.750 57.280 60.920 57.970 ;
        RECT 61.540 57.280 61.710 57.970 ;
        RECT 64.705 57.280 64.875 57.970 ;
        RECT 65.495 57.280 65.665 57.970 ;
        RECT 66.085 57.280 66.255 57.970 ;
        RECT 66.875 57.280 67.045 57.970 ;
        RECT 70.030 57.280 70.200 57.970 ;
        RECT 70.820 57.280 70.990 57.970 ;
        RECT 71.410 57.280 71.580 57.970 ;
        RECT 72.200 57.280 72.370 57.970 ;
        RECT 75.365 57.280 75.535 57.970 ;
        RECT 76.155 57.280 76.325 57.970 ;
        RECT 76.745 57.280 76.915 57.970 ;
        RECT 77.535 57.280 77.705 57.970 ;
        RECT 80.690 57.280 80.860 57.970 ;
        RECT 81.480 57.280 81.650 57.970 ;
        RECT 82.070 57.280 82.240 57.970 ;
        RECT 82.860 57.280 83.030 57.970 ;
        RECT 86.025 57.280 86.195 57.970 ;
        RECT 86.815 57.280 86.985 57.970 ;
        RECT 87.405 57.280 87.575 57.970 ;
        RECT 88.195 57.280 88.365 57.970 ;
        RECT 91.350 57.280 91.520 57.970 ;
        RECT 92.140 57.280 92.310 57.970 ;
        RECT 92.730 57.280 92.900 57.970 ;
        RECT 93.520 57.280 93.690 57.970 ;
        RECT 96.685 57.280 96.855 57.970 ;
        RECT 97.475 57.280 97.645 57.970 ;
        RECT 98.065 57.280 98.235 57.970 ;
        RECT 98.855 57.280 99.025 57.970 ;
        RECT 102.010 57.280 102.180 57.970 ;
        RECT 102.800 57.280 102.970 57.970 ;
        RECT 103.390 57.280 103.560 57.970 ;
        RECT 104.180 57.280 104.350 57.970 ;
        RECT 107.345 57.280 107.515 57.970 ;
        RECT 108.135 57.280 108.305 57.970 ;
        RECT 108.725 57.280 108.895 57.970 ;
        RECT 109.515 57.280 109.685 57.970 ;
        RECT 112.670 57.280 112.840 57.970 ;
        RECT 113.460 57.280 113.630 57.970 ;
        RECT 114.050 57.280 114.220 57.970 ;
        RECT 114.840 57.280 115.010 57.970 ;
        RECT 118.005 57.280 118.175 57.970 ;
        RECT 118.795 57.280 118.965 57.970 ;
        RECT 119.385 57.280 119.555 57.970 ;
        RECT 120.175 57.280 120.345 57.970 ;
        RECT 123.330 57.280 123.500 57.970 ;
        RECT 124.120 57.280 124.290 57.970 ;
        RECT 124.710 57.280 124.880 57.970 ;
        RECT 125.500 57.280 125.670 57.970 ;
        RECT 16.045 56.695 21.840 56.700 ;
        RECT 11.930 54.975 12.260 56.630 ;
        RECT 13.570 54.975 13.820 56.630 ;
        RECT 16.005 56.525 21.840 56.695 ;
        RECT 16.005 55.285 16.335 56.525 ;
        RECT 17.565 55.285 17.895 56.525 ;
        RECT 19.125 55.285 19.455 56.525 ;
        RECT 20.685 55.285 21.015 56.525 ;
        RECT 6.515 53.725 7.325 54.055 ;
        RECT 3.215 53.355 3.595 53.645 ;
        RECT 3.305 52.585 3.595 53.355 ;
        RECT 4.205 53.065 4.515 53.495 ;
        RECT 6.995 53.385 7.325 53.725 ;
        RECT 7.495 53.985 8.165 54.395 ;
        RECT 7.495 53.065 7.825 53.985 ;
        RECT 4.205 52.755 6.120 53.065 ;
        RECT 4.810 52.735 6.120 52.755 ;
        RECT 6.290 52.735 9.740 53.065 ;
        RECT 3.305 52.335 4.640 52.585 ;
        RECT 3.305 51.325 3.595 52.335 ;
        RECT 4.810 52.165 5.140 52.735 ;
        RECT 4.205 51.835 5.140 52.165 ;
        RECT 4.205 51.325 4.515 51.835 ;
        RECT 6.290 51.185 6.620 52.735 ;
        RECT 7.850 51.185 8.180 52.735 ;
        RECT 9.410 51.105 9.740 52.735 ;
        RECT 11.015 52.140 11.960 52.470 ;
        RECT 12.130 52.370 12.380 54.345 ;
        RECT 14.565 52.795 14.895 54.035 ;
        RECT 16.125 52.795 16.455 54.035 ;
        RECT 17.685 52.795 18.015 54.035 ;
        RECT 19.245 52.795 19.575 54.035 ;
        RECT 14.565 52.625 20.400 52.795 ;
        RECT 16.175 52.610 20.400 52.625 ;
        RECT 14.645 52.405 15.945 52.435 ;
        RECT 12.130 52.200 12.685 52.370 ;
        RECT 12.455 51.960 12.685 52.200 ;
        RECT 13.600 52.170 20.050 52.405 ;
        RECT 12.090 51.130 12.685 51.960 ;
        RECT 14.485 51.985 19.515 51.990 ;
        RECT 20.230 51.985 20.400 52.610 ;
        RECT 31.475 52.490 32.185 57.065 ;
        RECT 32.725 55.485 32.895 56.525 ;
        RECT 33.515 55.485 33.685 56.525 ;
        RECT 34.105 55.485 34.275 56.525 ;
        RECT 34.895 55.485 35.065 56.525 ;
        RECT 32.725 52.930 32.895 53.970 ;
        RECT 33.515 52.930 33.685 53.970 ;
        RECT 34.105 52.930 34.275 53.970 ;
        RECT 34.895 52.930 35.065 53.970 ;
        RECT 35.610 52.490 36.320 57.065 ;
        RECT 36.800 52.475 37.510 57.050 ;
        RECT 38.050 55.485 38.220 56.525 ;
        RECT 38.840 55.485 39.010 56.525 ;
        RECT 39.430 55.485 39.600 56.525 ;
        RECT 40.220 55.485 40.390 56.525 ;
        RECT 38.280 55.100 38.780 55.270 ;
        RECT 39.660 55.100 40.160 55.270 ;
        RECT 38.280 54.185 38.780 54.355 ;
        RECT 39.660 54.185 40.160 54.355 ;
        RECT 38.050 52.930 38.220 53.970 ;
        RECT 38.840 52.930 39.010 53.970 ;
        RECT 39.430 52.930 39.600 53.970 ;
        RECT 40.220 52.930 40.390 53.970 ;
        RECT 40.935 52.470 41.645 57.045 ;
        RECT 42.135 52.475 42.845 57.050 ;
        RECT 43.385 55.485 43.555 56.525 ;
        RECT 44.175 55.485 44.345 56.525 ;
        RECT 44.765 55.485 44.935 56.525 ;
        RECT 45.555 55.485 45.725 56.525 ;
        RECT 43.615 55.100 44.115 55.270 ;
        RECT 44.995 55.100 45.495 55.270 ;
        RECT 43.615 54.185 44.115 54.355 ;
        RECT 44.995 54.185 45.495 54.355 ;
        RECT 43.385 52.930 43.555 53.970 ;
        RECT 44.175 52.930 44.345 53.970 ;
        RECT 44.765 52.930 44.935 53.970 ;
        RECT 45.555 52.930 45.725 53.970 ;
        RECT 46.270 52.470 46.980 57.045 ;
        RECT 47.460 52.475 48.170 57.050 ;
        RECT 48.710 55.485 48.880 56.525 ;
        RECT 49.500 55.485 49.670 56.525 ;
        RECT 50.090 55.485 50.260 56.525 ;
        RECT 50.880 55.485 51.050 56.525 ;
        RECT 48.940 55.100 49.440 55.270 ;
        RECT 50.320 55.100 50.820 55.270 ;
        RECT 48.940 54.185 49.440 54.355 ;
        RECT 50.320 54.185 50.820 54.355 ;
        RECT 48.710 52.930 48.880 53.970 ;
        RECT 49.500 52.930 49.670 53.970 ;
        RECT 50.090 52.930 50.260 53.970 ;
        RECT 50.880 52.930 51.050 53.970 ;
        RECT 51.595 52.470 52.305 57.045 ;
        RECT 52.795 52.475 53.505 57.050 ;
        RECT 54.045 55.485 54.215 56.525 ;
        RECT 54.835 55.485 55.005 56.525 ;
        RECT 55.425 55.485 55.595 56.525 ;
        RECT 56.215 55.485 56.385 56.525 ;
        RECT 54.275 55.100 54.775 55.270 ;
        RECT 55.655 55.100 56.155 55.270 ;
        RECT 54.275 54.185 54.775 54.355 ;
        RECT 55.655 54.185 56.155 54.355 ;
        RECT 54.045 52.930 54.215 53.970 ;
        RECT 54.835 52.930 55.005 53.970 ;
        RECT 55.425 52.930 55.595 53.970 ;
        RECT 56.215 52.930 56.385 53.970 ;
        RECT 56.930 52.470 57.640 57.045 ;
        RECT 58.120 52.475 58.830 57.050 ;
        RECT 59.370 55.485 59.540 56.525 ;
        RECT 60.160 55.485 60.330 56.525 ;
        RECT 60.750 55.485 60.920 56.525 ;
        RECT 61.540 55.485 61.710 56.525 ;
        RECT 59.600 55.100 60.100 55.270 ;
        RECT 60.980 55.100 61.480 55.270 ;
        RECT 59.600 54.185 60.100 54.355 ;
        RECT 60.980 54.185 61.480 54.355 ;
        RECT 59.370 52.930 59.540 53.970 ;
        RECT 60.160 52.930 60.330 53.970 ;
        RECT 60.750 52.930 60.920 53.970 ;
        RECT 61.540 52.930 61.710 53.970 ;
        RECT 62.255 52.470 62.965 57.045 ;
        RECT 63.455 52.475 64.165 57.050 ;
        RECT 64.705 55.485 64.875 56.525 ;
        RECT 65.495 55.485 65.665 56.525 ;
        RECT 66.085 55.485 66.255 56.525 ;
        RECT 66.875 55.485 67.045 56.525 ;
        RECT 64.935 55.100 65.435 55.270 ;
        RECT 66.315 55.100 66.815 55.270 ;
        RECT 64.935 54.185 65.435 54.355 ;
        RECT 66.315 54.185 66.815 54.355 ;
        RECT 64.705 52.930 64.875 53.970 ;
        RECT 65.495 52.930 65.665 53.970 ;
        RECT 66.085 52.930 66.255 53.970 ;
        RECT 66.875 52.930 67.045 53.970 ;
        RECT 67.590 52.470 68.300 57.045 ;
        RECT 68.780 52.475 69.490 57.050 ;
        RECT 70.030 55.485 70.200 56.525 ;
        RECT 70.820 55.485 70.990 56.525 ;
        RECT 71.410 55.485 71.580 56.525 ;
        RECT 72.200 55.485 72.370 56.525 ;
        RECT 70.260 55.100 70.760 55.270 ;
        RECT 71.640 55.100 72.140 55.270 ;
        RECT 70.260 54.185 70.760 54.355 ;
        RECT 71.640 54.185 72.140 54.355 ;
        RECT 70.030 52.930 70.200 53.970 ;
        RECT 70.820 52.930 70.990 53.970 ;
        RECT 71.410 52.930 71.580 53.970 ;
        RECT 72.200 52.930 72.370 53.970 ;
        RECT 72.915 52.470 73.625 57.045 ;
        RECT 74.115 52.475 74.825 57.050 ;
        RECT 75.365 55.485 75.535 56.525 ;
        RECT 76.155 55.485 76.325 56.525 ;
        RECT 76.745 55.485 76.915 56.525 ;
        RECT 77.535 55.485 77.705 56.525 ;
        RECT 75.595 55.100 76.095 55.270 ;
        RECT 76.975 55.100 77.475 55.270 ;
        RECT 75.595 54.185 76.095 54.355 ;
        RECT 76.975 54.185 77.475 54.355 ;
        RECT 75.365 52.930 75.535 53.970 ;
        RECT 76.155 52.930 76.325 53.970 ;
        RECT 76.745 52.930 76.915 53.970 ;
        RECT 77.535 52.930 77.705 53.970 ;
        RECT 78.250 52.470 78.960 57.045 ;
        RECT 79.440 52.475 80.150 57.050 ;
        RECT 80.690 55.485 80.860 56.525 ;
        RECT 81.480 55.485 81.650 56.525 ;
        RECT 82.070 55.485 82.240 56.525 ;
        RECT 82.860 55.485 83.030 56.525 ;
        RECT 80.920 55.100 81.420 55.270 ;
        RECT 82.300 55.100 82.800 55.270 ;
        RECT 80.920 54.185 81.420 54.355 ;
        RECT 82.300 54.185 82.800 54.355 ;
        RECT 80.690 52.930 80.860 53.970 ;
        RECT 81.480 52.930 81.650 53.970 ;
        RECT 82.070 52.930 82.240 53.970 ;
        RECT 82.860 52.930 83.030 53.970 ;
        RECT 83.575 52.470 84.285 57.045 ;
        RECT 84.775 52.475 85.485 57.050 ;
        RECT 86.025 55.485 86.195 56.525 ;
        RECT 86.815 55.485 86.985 56.525 ;
        RECT 87.405 55.485 87.575 56.525 ;
        RECT 88.195 55.485 88.365 56.525 ;
        RECT 86.255 55.100 86.755 55.270 ;
        RECT 87.635 55.100 88.135 55.270 ;
        RECT 86.255 54.185 86.755 54.355 ;
        RECT 87.635 54.185 88.135 54.355 ;
        RECT 86.025 52.930 86.195 53.970 ;
        RECT 86.815 52.930 86.985 53.970 ;
        RECT 87.405 52.930 87.575 53.970 ;
        RECT 88.195 52.930 88.365 53.970 ;
        RECT 88.910 52.470 89.620 57.045 ;
        RECT 90.100 52.475 90.810 57.050 ;
        RECT 91.350 55.485 91.520 56.525 ;
        RECT 92.140 55.485 92.310 56.525 ;
        RECT 92.730 55.485 92.900 56.525 ;
        RECT 93.520 55.485 93.690 56.525 ;
        RECT 91.580 55.100 92.080 55.270 ;
        RECT 92.960 55.100 93.460 55.270 ;
        RECT 91.580 54.185 92.080 54.355 ;
        RECT 92.960 54.185 93.460 54.355 ;
        RECT 91.350 52.930 91.520 53.970 ;
        RECT 92.140 52.930 92.310 53.970 ;
        RECT 92.730 52.930 92.900 53.970 ;
        RECT 93.520 52.930 93.690 53.970 ;
        RECT 94.235 52.470 94.945 57.045 ;
        RECT 95.435 52.475 96.145 57.050 ;
        RECT 96.685 55.485 96.855 56.525 ;
        RECT 97.475 55.485 97.645 56.525 ;
        RECT 98.065 55.485 98.235 56.525 ;
        RECT 98.855 55.485 99.025 56.525 ;
        RECT 96.915 55.100 97.415 55.270 ;
        RECT 98.295 55.100 98.795 55.270 ;
        RECT 96.915 54.185 97.415 54.355 ;
        RECT 98.295 54.185 98.795 54.355 ;
        RECT 96.685 52.930 96.855 53.970 ;
        RECT 97.475 52.930 97.645 53.970 ;
        RECT 98.065 52.930 98.235 53.970 ;
        RECT 98.855 52.930 99.025 53.970 ;
        RECT 99.570 52.470 100.280 57.045 ;
        RECT 100.760 52.475 101.470 57.050 ;
        RECT 102.010 55.485 102.180 56.525 ;
        RECT 102.800 55.485 102.970 56.525 ;
        RECT 103.390 55.485 103.560 56.525 ;
        RECT 104.180 55.485 104.350 56.525 ;
        RECT 102.240 55.100 102.740 55.270 ;
        RECT 103.620 55.100 104.120 55.270 ;
        RECT 102.240 54.185 102.740 54.355 ;
        RECT 103.620 54.185 104.120 54.355 ;
        RECT 102.010 52.930 102.180 53.970 ;
        RECT 102.800 52.930 102.970 53.970 ;
        RECT 103.390 52.930 103.560 53.970 ;
        RECT 104.180 52.930 104.350 53.970 ;
        RECT 104.895 52.470 105.605 57.045 ;
        RECT 106.095 52.475 106.805 57.050 ;
        RECT 107.345 55.485 107.515 56.525 ;
        RECT 108.135 55.485 108.305 56.525 ;
        RECT 108.725 55.485 108.895 56.525 ;
        RECT 109.515 55.485 109.685 56.525 ;
        RECT 107.575 55.100 108.075 55.270 ;
        RECT 108.955 55.100 109.455 55.270 ;
        RECT 107.575 54.185 108.075 54.355 ;
        RECT 108.955 54.185 109.455 54.355 ;
        RECT 107.345 52.930 107.515 53.970 ;
        RECT 108.135 52.930 108.305 53.970 ;
        RECT 108.725 52.930 108.895 53.970 ;
        RECT 109.515 52.930 109.685 53.970 ;
        RECT 110.230 52.470 110.940 57.045 ;
        RECT 111.420 52.475 112.130 57.050 ;
        RECT 112.670 55.485 112.840 56.525 ;
        RECT 113.460 55.485 113.630 56.525 ;
        RECT 114.050 55.485 114.220 56.525 ;
        RECT 114.840 55.485 115.010 56.525 ;
        RECT 112.900 55.100 113.400 55.270 ;
        RECT 114.280 55.100 114.780 55.270 ;
        RECT 112.900 54.185 113.400 54.355 ;
        RECT 114.280 54.185 114.780 54.355 ;
        RECT 112.670 52.930 112.840 53.970 ;
        RECT 113.460 52.930 113.630 53.970 ;
        RECT 114.050 52.930 114.220 53.970 ;
        RECT 114.840 52.930 115.010 53.970 ;
        RECT 115.555 52.470 116.265 57.045 ;
        RECT 116.755 52.475 117.465 57.050 ;
        RECT 118.005 55.485 118.175 56.525 ;
        RECT 118.795 55.485 118.965 56.525 ;
        RECT 119.385 55.485 119.555 56.525 ;
        RECT 120.175 55.485 120.345 56.525 ;
        RECT 118.235 55.100 118.735 55.270 ;
        RECT 119.615 55.100 120.115 55.270 ;
        RECT 118.235 54.185 118.735 54.355 ;
        RECT 119.615 54.185 120.115 54.355 ;
        RECT 118.005 52.930 118.175 53.970 ;
        RECT 118.795 52.930 118.965 53.970 ;
        RECT 119.385 52.930 119.555 53.970 ;
        RECT 120.175 52.930 120.345 53.970 ;
        RECT 120.890 52.470 121.600 57.045 ;
        RECT 122.080 52.490 122.790 57.065 ;
        RECT 123.330 55.485 123.500 56.525 ;
        RECT 124.120 55.485 124.290 56.525 ;
        RECT 124.710 55.485 124.880 56.525 ;
        RECT 125.500 55.485 125.670 56.525 ;
        RECT 123.330 52.930 123.500 53.970 ;
        RECT 124.120 52.930 124.290 53.970 ;
        RECT 124.710 52.930 124.880 53.970 ;
        RECT 125.500 52.930 125.670 53.970 ;
        RECT 126.215 52.490 126.925 57.065 ;
        RECT 14.485 51.820 20.400 51.985 ;
        RECT 14.485 51.320 14.695 51.820 ;
        RECT 16.045 51.815 20.400 51.820 ;
        RECT 16.045 51.805 20.260 51.815 ;
        RECT 16.045 51.320 16.255 51.805 ;
        RECT 17.605 51.320 17.815 51.805 ;
        RECT 19.205 51.320 19.855 51.805 ;
        RECT 32.725 51.485 32.895 52.175 ;
        RECT 33.515 51.485 33.685 52.175 ;
        RECT 34.105 51.485 34.275 52.175 ;
        RECT 34.895 51.485 35.065 52.175 ;
        RECT 38.050 51.485 38.220 52.175 ;
        RECT 38.840 51.485 39.010 52.175 ;
        RECT 39.430 51.485 39.600 52.175 ;
        RECT 40.220 51.485 40.390 52.175 ;
        RECT 43.385 51.485 43.555 52.175 ;
        RECT 44.175 51.485 44.345 52.175 ;
        RECT 44.765 51.485 44.935 52.175 ;
        RECT 45.555 51.485 45.725 52.175 ;
        RECT 48.710 51.485 48.880 52.175 ;
        RECT 49.500 51.485 49.670 52.175 ;
        RECT 50.090 51.485 50.260 52.175 ;
        RECT 50.880 51.485 51.050 52.175 ;
        RECT 54.045 51.485 54.215 52.175 ;
        RECT 54.835 51.485 55.005 52.175 ;
        RECT 55.425 51.485 55.595 52.175 ;
        RECT 56.215 51.485 56.385 52.175 ;
        RECT 59.370 51.485 59.540 52.175 ;
        RECT 60.160 51.485 60.330 52.175 ;
        RECT 60.750 51.485 60.920 52.175 ;
        RECT 61.540 51.485 61.710 52.175 ;
        RECT 64.705 51.485 64.875 52.175 ;
        RECT 65.495 51.485 65.665 52.175 ;
        RECT 66.085 51.485 66.255 52.175 ;
        RECT 66.875 51.485 67.045 52.175 ;
        RECT 70.030 51.485 70.200 52.175 ;
        RECT 70.820 51.485 70.990 52.175 ;
        RECT 71.410 51.485 71.580 52.175 ;
        RECT 72.200 51.485 72.370 52.175 ;
        RECT 75.365 51.485 75.535 52.175 ;
        RECT 76.155 51.485 76.325 52.175 ;
        RECT 76.745 51.485 76.915 52.175 ;
        RECT 77.535 51.485 77.705 52.175 ;
        RECT 80.690 51.485 80.860 52.175 ;
        RECT 81.480 51.485 81.650 52.175 ;
        RECT 82.070 51.485 82.240 52.175 ;
        RECT 82.860 51.485 83.030 52.175 ;
        RECT 86.025 51.485 86.195 52.175 ;
        RECT 86.815 51.485 86.985 52.175 ;
        RECT 87.405 51.485 87.575 52.175 ;
        RECT 88.195 51.485 88.365 52.175 ;
        RECT 91.350 51.485 91.520 52.175 ;
        RECT 92.140 51.485 92.310 52.175 ;
        RECT 92.730 51.485 92.900 52.175 ;
        RECT 93.520 51.485 93.690 52.175 ;
        RECT 96.685 51.485 96.855 52.175 ;
        RECT 97.475 51.485 97.645 52.175 ;
        RECT 98.065 51.485 98.235 52.175 ;
        RECT 98.855 51.485 99.025 52.175 ;
        RECT 102.010 51.485 102.180 52.175 ;
        RECT 102.800 51.485 102.970 52.175 ;
        RECT 103.390 51.485 103.560 52.175 ;
        RECT 104.180 51.485 104.350 52.175 ;
        RECT 107.345 51.485 107.515 52.175 ;
        RECT 108.135 51.485 108.305 52.175 ;
        RECT 108.725 51.485 108.895 52.175 ;
        RECT 109.515 51.485 109.685 52.175 ;
        RECT 112.670 51.485 112.840 52.175 ;
        RECT 113.460 51.485 113.630 52.175 ;
        RECT 114.050 51.485 114.220 52.175 ;
        RECT 114.840 51.485 115.010 52.175 ;
        RECT 118.005 51.485 118.175 52.175 ;
        RECT 118.795 51.485 118.965 52.175 ;
        RECT 119.385 51.485 119.555 52.175 ;
        RECT 120.175 51.485 120.345 52.175 ;
        RECT 123.330 51.485 123.500 52.175 ;
        RECT 124.120 51.485 124.290 52.175 ;
        RECT 124.710 51.485 124.880 52.175 ;
        RECT 125.500 51.485 125.670 52.175 ;
        RECT 38.280 51.145 38.780 51.315 ;
        RECT 39.660 51.145 40.160 51.315 ;
        RECT 43.615 51.145 44.115 51.315 ;
        RECT 44.995 51.145 45.495 51.315 ;
        RECT 48.940 51.145 49.440 51.315 ;
        RECT 50.320 51.145 50.820 51.315 ;
        RECT 54.275 51.145 54.775 51.315 ;
        RECT 55.655 51.145 56.155 51.315 ;
        RECT 59.600 51.145 60.100 51.315 ;
        RECT 60.980 51.145 61.480 51.315 ;
        RECT 64.935 51.145 65.435 51.315 ;
        RECT 66.315 51.145 66.815 51.315 ;
        RECT 70.260 51.145 70.760 51.315 ;
        RECT 71.640 51.145 72.140 51.315 ;
        RECT 75.595 51.145 76.095 51.315 ;
        RECT 76.975 51.145 77.475 51.315 ;
        RECT 80.920 51.145 81.420 51.315 ;
        RECT 82.300 51.145 82.800 51.315 ;
        RECT 86.255 51.145 86.755 51.315 ;
        RECT 87.635 51.145 88.135 51.315 ;
        RECT 91.580 51.145 92.080 51.315 ;
        RECT 92.960 51.145 93.460 51.315 ;
        RECT 96.915 51.145 97.415 51.315 ;
        RECT 98.295 51.145 98.795 51.315 ;
        RECT 102.240 51.145 102.740 51.315 ;
        RECT 103.620 51.145 104.120 51.315 ;
        RECT 107.575 51.145 108.075 51.315 ;
        RECT 108.955 51.145 109.455 51.315 ;
        RECT 112.900 51.145 113.400 51.315 ;
        RECT 114.280 51.145 114.780 51.315 ;
        RECT 118.235 51.145 118.735 51.315 ;
        RECT 119.615 51.145 120.115 51.315 ;
        RECT 38.280 50.605 38.780 50.775 ;
        RECT 39.660 50.605 40.160 50.775 ;
        RECT 43.615 50.605 44.115 50.775 ;
        RECT 44.995 50.605 45.495 50.775 ;
        RECT 48.940 50.605 49.440 50.775 ;
        RECT 50.320 50.605 50.820 50.775 ;
        RECT 54.275 50.605 54.775 50.775 ;
        RECT 55.655 50.605 56.155 50.775 ;
        RECT 59.600 50.605 60.100 50.775 ;
        RECT 60.980 50.605 61.480 50.775 ;
        RECT 64.935 50.605 65.435 50.775 ;
        RECT 66.315 50.605 66.815 50.775 ;
        RECT 70.260 50.605 70.760 50.775 ;
        RECT 71.640 50.605 72.140 50.775 ;
        RECT 75.595 50.605 76.095 50.775 ;
        RECT 76.975 50.605 77.475 50.775 ;
        RECT 80.920 50.605 81.420 50.775 ;
        RECT 82.300 50.605 82.800 50.775 ;
        RECT 86.255 50.605 86.755 50.775 ;
        RECT 87.635 50.605 88.135 50.775 ;
        RECT 91.580 50.605 92.080 50.775 ;
        RECT 92.960 50.605 93.460 50.775 ;
        RECT 96.915 50.605 97.415 50.775 ;
        RECT 98.295 50.605 98.795 50.775 ;
        RECT 102.240 50.605 102.740 50.775 ;
        RECT 103.620 50.605 104.120 50.775 ;
        RECT 107.575 50.605 108.075 50.775 ;
        RECT 108.955 50.605 109.455 50.775 ;
        RECT 112.900 50.605 113.400 50.775 ;
        RECT 114.280 50.605 114.780 50.775 ;
        RECT 118.235 50.605 118.735 50.775 ;
        RECT 119.615 50.605 120.115 50.775 ;
        RECT 2.825 48.445 3.155 49.995 ;
        RECT 4.385 48.445 4.715 49.995 ;
        RECT 5.945 48.445 6.275 50.075 ;
        RECT 8.845 49.005 9.175 50.075 ;
        RECT 10.450 49.175 10.780 50.075 ;
        RECT 11.930 49.360 12.180 50.095 ;
        RECT 13.490 49.360 14.075 50.095 ;
        RECT 11.930 49.190 14.075 49.360 ;
        RECT 15.925 49.365 16.135 49.860 ;
        RECT 17.485 49.365 17.695 49.860 ;
        RECT 19.045 49.365 19.255 49.860 ;
        RECT 20.645 49.365 21.295 49.860 ;
        RECT 32.725 49.745 32.895 50.435 ;
        RECT 33.515 49.745 33.685 50.435 ;
        RECT 34.105 49.745 34.275 50.435 ;
        RECT 34.895 49.745 35.065 50.435 ;
        RECT 38.050 49.745 38.220 50.435 ;
        RECT 38.840 49.745 39.010 50.435 ;
        RECT 39.430 49.745 39.600 50.435 ;
        RECT 40.220 49.745 40.390 50.435 ;
        RECT 43.385 49.745 43.555 50.435 ;
        RECT 44.175 49.745 44.345 50.435 ;
        RECT 44.765 49.745 44.935 50.435 ;
        RECT 45.555 49.745 45.725 50.435 ;
        RECT 48.710 49.745 48.880 50.435 ;
        RECT 49.500 49.745 49.670 50.435 ;
        RECT 50.090 49.745 50.260 50.435 ;
        RECT 50.880 49.745 51.050 50.435 ;
        RECT 54.045 49.745 54.215 50.435 ;
        RECT 54.835 49.745 55.005 50.435 ;
        RECT 55.425 49.745 55.595 50.435 ;
        RECT 56.215 49.745 56.385 50.435 ;
        RECT 59.370 49.745 59.540 50.435 ;
        RECT 60.160 49.745 60.330 50.435 ;
        RECT 60.750 49.745 60.920 50.435 ;
        RECT 61.540 49.745 61.710 50.435 ;
        RECT 64.705 49.745 64.875 50.435 ;
        RECT 65.495 49.745 65.665 50.435 ;
        RECT 66.085 49.745 66.255 50.435 ;
        RECT 66.875 49.745 67.045 50.435 ;
        RECT 70.030 49.745 70.200 50.435 ;
        RECT 70.820 49.745 70.990 50.435 ;
        RECT 71.410 49.745 71.580 50.435 ;
        RECT 72.200 49.745 72.370 50.435 ;
        RECT 75.365 49.745 75.535 50.435 ;
        RECT 76.155 49.745 76.325 50.435 ;
        RECT 76.745 49.745 76.915 50.435 ;
        RECT 77.535 49.745 77.705 50.435 ;
        RECT 80.690 49.745 80.860 50.435 ;
        RECT 81.480 49.745 81.650 50.435 ;
        RECT 82.070 49.745 82.240 50.435 ;
        RECT 82.860 49.745 83.030 50.435 ;
        RECT 86.025 49.745 86.195 50.435 ;
        RECT 86.815 49.745 86.985 50.435 ;
        RECT 87.405 49.745 87.575 50.435 ;
        RECT 88.195 49.745 88.365 50.435 ;
        RECT 91.350 49.745 91.520 50.435 ;
        RECT 92.140 49.745 92.310 50.435 ;
        RECT 92.730 49.745 92.900 50.435 ;
        RECT 93.520 49.745 93.690 50.435 ;
        RECT 96.685 49.745 96.855 50.435 ;
        RECT 97.475 49.745 97.645 50.435 ;
        RECT 98.065 49.745 98.235 50.435 ;
        RECT 98.855 49.745 99.025 50.435 ;
        RECT 102.010 49.745 102.180 50.435 ;
        RECT 102.800 49.745 102.970 50.435 ;
        RECT 103.390 49.745 103.560 50.435 ;
        RECT 104.180 49.745 104.350 50.435 ;
        RECT 107.345 49.745 107.515 50.435 ;
        RECT 108.135 49.745 108.305 50.435 ;
        RECT 108.725 49.745 108.895 50.435 ;
        RECT 109.515 49.745 109.685 50.435 ;
        RECT 112.670 49.745 112.840 50.435 ;
        RECT 113.460 49.745 113.630 50.435 ;
        RECT 114.050 49.745 114.220 50.435 ;
        RECT 114.840 49.745 115.010 50.435 ;
        RECT 118.005 49.745 118.175 50.435 ;
        RECT 118.795 49.745 118.965 50.435 ;
        RECT 119.385 49.745 119.555 50.435 ;
        RECT 120.175 49.745 120.345 50.435 ;
        RECT 123.330 49.745 123.500 50.435 ;
        RECT 124.120 49.745 124.290 50.435 ;
        RECT 124.710 49.745 124.880 50.435 ;
        RECT 125.500 49.745 125.670 50.435 ;
        RECT 15.925 49.190 21.840 49.365 ;
        RECT 7.990 48.445 8.320 49.005 ;
        RECT 2.825 48.115 8.320 48.445 ;
        RECT 3.215 45.505 3.505 47.945 ;
        RECT 6.515 45.915 6.845 48.115 ;
        RECT 7.990 47.655 8.320 48.115 ;
        RECT 8.845 48.675 10.370 49.005 ;
        RECT 7.015 46.920 7.825 47.250 ;
        RECT 7.495 46.255 7.825 46.920 ;
        RECT 8.845 46.855 9.175 48.675 ;
        RECT 10.540 48.505 10.780 49.175 ;
        RECT 13.905 49.040 14.075 49.190 ;
        RECT 13.905 49.010 14.605 49.040 ;
        RECT 11.015 48.840 13.725 49.010 ;
        RECT 13.905 48.775 21.490 49.010 ;
        RECT 13.905 48.660 15.710 48.775 ;
        RECT 10.450 46.855 10.780 48.505 ;
        RECT 11.930 48.490 15.710 48.660 ;
        RECT 21.670 48.560 21.840 49.190 ;
        RECT 16.045 48.555 21.840 48.560 ;
        RECT 11.930 46.835 12.260 48.490 ;
        RECT 13.570 46.835 13.820 48.490 ;
        RECT 16.005 48.385 21.840 48.555 ;
        RECT 16.005 47.145 16.335 48.385 ;
        RECT 17.565 47.145 17.895 48.385 ;
        RECT 19.125 47.145 19.455 48.385 ;
        RECT 20.685 47.145 21.015 48.385 ;
        RECT 6.515 45.585 7.325 45.915 ;
        RECT 3.215 45.215 3.595 45.505 ;
        RECT 3.305 44.445 3.595 45.215 ;
        RECT 4.205 44.925 4.515 45.355 ;
        RECT 6.995 45.245 7.325 45.585 ;
        RECT 7.495 45.845 8.165 46.255 ;
        RECT 7.495 44.925 7.825 45.845 ;
        RECT 4.205 44.615 6.120 44.925 ;
        RECT 4.810 44.595 6.120 44.615 ;
        RECT 6.290 44.595 9.740 44.925 ;
        RECT 3.305 44.195 4.640 44.445 ;
        RECT 3.305 43.185 3.595 44.195 ;
        RECT 4.810 44.025 5.140 44.595 ;
        RECT 4.205 43.695 5.140 44.025 ;
        RECT 4.205 43.185 4.515 43.695 ;
        RECT 6.290 43.045 6.620 44.595 ;
        RECT 7.850 43.045 8.180 44.595 ;
        RECT 9.410 42.965 9.740 44.595 ;
        RECT 11.015 44.000 11.960 44.330 ;
        RECT 12.130 44.230 12.380 46.205 ;
        RECT 14.565 44.655 14.895 45.895 ;
        RECT 16.125 44.655 16.455 45.895 ;
        RECT 17.685 44.655 18.015 45.895 ;
        RECT 19.245 44.655 19.575 45.895 ;
        RECT 31.475 44.955 32.185 49.530 ;
        RECT 32.725 47.950 32.895 48.990 ;
        RECT 33.515 47.950 33.685 48.990 ;
        RECT 34.105 47.950 34.275 48.990 ;
        RECT 34.895 47.950 35.065 48.990 ;
        RECT 32.725 45.395 32.895 46.435 ;
        RECT 33.515 45.395 33.685 46.435 ;
        RECT 34.105 45.395 34.275 46.435 ;
        RECT 34.895 45.395 35.065 46.435 ;
        RECT 35.610 44.955 36.320 49.530 ;
        RECT 36.800 44.940 37.510 49.515 ;
        RECT 38.050 47.950 38.220 48.990 ;
        RECT 38.840 47.950 39.010 48.990 ;
        RECT 39.430 47.950 39.600 48.990 ;
        RECT 40.220 47.950 40.390 48.990 ;
        RECT 38.280 47.565 38.780 47.735 ;
        RECT 39.660 47.565 40.160 47.735 ;
        RECT 38.280 46.650 38.780 46.820 ;
        RECT 39.660 46.650 40.160 46.820 ;
        RECT 38.050 45.395 38.220 46.435 ;
        RECT 38.840 45.395 39.010 46.435 ;
        RECT 39.430 45.395 39.600 46.435 ;
        RECT 40.220 45.395 40.390 46.435 ;
        RECT 40.935 44.935 41.645 49.510 ;
        RECT 42.135 44.940 42.845 49.515 ;
        RECT 43.385 47.950 43.555 48.990 ;
        RECT 44.175 47.950 44.345 48.990 ;
        RECT 44.765 47.950 44.935 48.990 ;
        RECT 45.555 47.950 45.725 48.990 ;
        RECT 43.615 47.565 44.115 47.735 ;
        RECT 44.995 47.565 45.495 47.735 ;
        RECT 43.615 46.650 44.115 46.820 ;
        RECT 44.995 46.650 45.495 46.820 ;
        RECT 43.385 45.395 43.555 46.435 ;
        RECT 44.175 45.395 44.345 46.435 ;
        RECT 44.765 45.395 44.935 46.435 ;
        RECT 45.555 45.395 45.725 46.435 ;
        RECT 46.270 44.935 46.980 49.510 ;
        RECT 47.460 44.940 48.170 49.515 ;
        RECT 48.710 47.950 48.880 48.990 ;
        RECT 49.500 47.950 49.670 48.990 ;
        RECT 50.090 47.950 50.260 48.990 ;
        RECT 50.880 47.950 51.050 48.990 ;
        RECT 48.940 47.565 49.440 47.735 ;
        RECT 50.320 47.565 50.820 47.735 ;
        RECT 48.940 46.650 49.440 46.820 ;
        RECT 50.320 46.650 50.820 46.820 ;
        RECT 48.710 45.395 48.880 46.435 ;
        RECT 49.500 45.395 49.670 46.435 ;
        RECT 50.090 45.395 50.260 46.435 ;
        RECT 50.880 45.395 51.050 46.435 ;
        RECT 51.595 44.935 52.305 49.510 ;
        RECT 52.795 44.940 53.505 49.515 ;
        RECT 54.045 47.950 54.215 48.990 ;
        RECT 54.835 47.950 55.005 48.990 ;
        RECT 55.425 47.950 55.595 48.990 ;
        RECT 56.215 47.950 56.385 48.990 ;
        RECT 54.275 47.565 54.775 47.735 ;
        RECT 55.655 47.565 56.155 47.735 ;
        RECT 54.275 46.650 54.775 46.820 ;
        RECT 55.655 46.650 56.155 46.820 ;
        RECT 54.045 45.395 54.215 46.435 ;
        RECT 54.835 45.395 55.005 46.435 ;
        RECT 55.425 45.395 55.595 46.435 ;
        RECT 56.215 45.395 56.385 46.435 ;
        RECT 56.930 44.935 57.640 49.510 ;
        RECT 58.120 44.940 58.830 49.515 ;
        RECT 59.370 47.950 59.540 48.990 ;
        RECT 60.160 47.950 60.330 48.990 ;
        RECT 60.750 47.950 60.920 48.990 ;
        RECT 61.540 47.950 61.710 48.990 ;
        RECT 59.600 47.565 60.100 47.735 ;
        RECT 60.980 47.565 61.480 47.735 ;
        RECT 59.600 46.650 60.100 46.820 ;
        RECT 60.980 46.650 61.480 46.820 ;
        RECT 59.370 45.395 59.540 46.435 ;
        RECT 60.160 45.395 60.330 46.435 ;
        RECT 60.750 45.395 60.920 46.435 ;
        RECT 61.540 45.395 61.710 46.435 ;
        RECT 62.255 44.935 62.965 49.510 ;
        RECT 63.455 44.940 64.165 49.515 ;
        RECT 64.705 47.950 64.875 48.990 ;
        RECT 65.495 47.950 65.665 48.990 ;
        RECT 66.085 47.950 66.255 48.990 ;
        RECT 66.875 47.950 67.045 48.990 ;
        RECT 64.935 47.565 65.435 47.735 ;
        RECT 66.315 47.565 66.815 47.735 ;
        RECT 64.935 46.650 65.435 46.820 ;
        RECT 66.315 46.650 66.815 46.820 ;
        RECT 64.705 45.395 64.875 46.435 ;
        RECT 65.495 45.395 65.665 46.435 ;
        RECT 66.085 45.395 66.255 46.435 ;
        RECT 66.875 45.395 67.045 46.435 ;
        RECT 67.590 44.935 68.300 49.510 ;
        RECT 68.780 44.940 69.490 49.515 ;
        RECT 70.030 47.950 70.200 48.990 ;
        RECT 70.820 47.950 70.990 48.990 ;
        RECT 71.410 47.950 71.580 48.990 ;
        RECT 72.200 47.950 72.370 48.990 ;
        RECT 70.260 47.565 70.760 47.735 ;
        RECT 71.640 47.565 72.140 47.735 ;
        RECT 70.260 46.650 70.760 46.820 ;
        RECT 71.640 46.650 72.140 46.820 ;
        RECT 70.030 45.395 70.200 46.435 ;
        RECT 70.820 45.395 70.990 46.435 ;
        RECT 71.410 45.395 71.580 46.435 ;
        RECT 72.200 45.395 72.370 46.435 ;
        RECT 72.915 44.935 73.625 49.510 ;
        RECT 74.115 44.940 74.825 49.515 ;
        RECT 75.365 47.950 75.535 48.990 ;
        RECT 76.155 47.950 76.325 48.990 ;
        RECT 76.745 47.950 76.915 48.990 ;
        RECT 77.535 47.950 77.705 48.990 ;
        RECT 75.595 47.565 76.095 47.735 ;
        RECT 76.975 47.565 77.475 47.735 ;
        RECT 75.595 46.650 76.095 46.820 ;
        RECT 76.975 46.650 77.475 46.820 ;
        RECT 75.365 45.395 75.535 46.435 ;
        RECT 76.155 45.395 76.325 46.435 ;
        RECT 76.745 45.395 76.915 46.435 ;
        RECT 77.535 45.395 77.705 46.435 ;
        RECT 78.250 44.935 78.960 49.510 ;
        RECT 79.440 44.940 80.150 49.515 ;
        RECT 80.690 47.950 80.860 48.990 ;
        RECT 81.480 47.950 81.650 48.990 ;
        RECT 82.070 47.950 82.240 48.990 ;
        RECT 82.860 47.950 83.030 48.990 ;
        RECT 80.920 47.565 81.420 47.735 ;
        RECT 82.300 47.565 82.800 47.735 ;
        RECT 80.920 46.650 81.420 46.820 ;
        RECT 82.300 46.650 82.800 46.820 ;
        RECT 80.690 45.395 80.860 46.435 ;
        RECT 81.480 45.395 81.650 46.435 ;
        RECT 82.070 45.395 82.240 46.435 ;
        RECT 82.860 45.395 83.030 46.435 ;
        RECT 83.575 44.935 84.285 49.510 ;
        RECT 84.775 44.940 85.485 49.515 ;
        RECT 86.025 47.950 86.195 48.990 ;
        RECT 86.815 47.950 86.985 48.990 ;
        RECT 87.405 47.950 87.575 48.990 ;
        RECT 88.195 47.950 88.365 48.990 ;
        RECT 86.255 47.565 86.755 47.735 ;
        RECT 87.635 47.565 88.135 47.735 ;
        RECT 86.255 46.650 86.755 46.820 ;
        RECT 87.635 46.650 88.135 46.820 ;
        RECT 86.025 45.395 86.195 46.435 ;
        RECT 86.815 45.395 86.985 46.435 ;
        RECT 87.405 45.395 87.575 46.435 ;
        RECT 88.195 45.395 88.365 46.435 ;
        RECT 88.910 44.935 89.620 49.510 ;
        RECT 90.100 44.940 90.810 49.515 ;
        RECT 91.350 47.950 91.520 48.990 ;
        RECT 92.140 47.950 92.310 48.990 ;
        RECT 92.730 47.950 92.900 48.990 ;
        RECT 93.520 47.950 93.690 48.990 ;
        RECT 91.580 47.565 92.080 47.735 ;
        RECT 92.960 47.565 93.460 47.735 ;
        RECT 91.580 46.650 92.080 46.820 ;
        RECT 92.960 46.650 93.460 46.820 ;
        RECT 91.350 45.395 91.520 46.435 ;
        RECT 92.140 45.395 92.310 46.435 ;
        RECT 92.730 45.395 92.900 46.435 ;
        RECT 93.520 45.395 93.690 46.435 ;
        RECT 94.235 44.935 94.945 49.510 ;
        RECT 95.435 44.940 96.145 49.515 ;
        RECT 96.685 47.950 96.855 48.990 ;
        RECT 97.475 47.950 97.645 48.990 ;
        RECT 98.065 47.950 98.235 48.990 ;
        RECT 98.855 47.950 99.025 48.990 ;
        RECT 96.915 47.565 97.415 47.735 ;
        RECT 98.295 47.565 98.795 47.735 ;
        RECT 96.915 46.650 97.415 46.820 ;
        RECT 98.295 46.650 98.795 46.820 ;
        RECT 96.685 45.395 96.855 46.435 ;
        RECT 97.475 45.395 97.645 46.435 ;
        RECT 98.065 45.395 98.235 46.435 ;
        RECT 98.855 45.395 99.025 46.435 ;
        RECT 99.570 44.935 100.280 49.510 ;
        RECT 100.760 44.940 101.470 49.515 ;
        RECT 102.010 47.950 102.180 48.990 ;
        RECT 102.800 47.950 102.970 48.990 ;
        RECT 103.390 47.950 103.560 48.990 ;
        RECT 104.180 47.950 104.350 48.990 ;
        RECT 102.240 47.565 102.740 47.735 ;
        RECT 103.620 47.565 104.120 47.735 ;
        RECT 102.240 46.650 102.740 46.820 ;
        RECT 103.620 46.650 104.120 46.820 ;
        RECT 102.010 45.395 102.180 46.435 ;
        RECT 102.800 45.395 102.970 46.435 ;
        RECT 103.390 45.395 103.560 46.435 ;
        RECT 104.180 45.395 104.350 46.435 ;
        RECT 104.895 44.935 105.605 49.510 ;
        RECT 106.095 44.940 106.805 49.515 ;
        RECT 107.345 47.950 107.515 48.990 ;
        RECT 108.135 47.950 108.305 48.990 ;
        RECT 108.725 47.950 108.895 48.990 ;
        RECT 109.515 47.950 109.685 48.990 ;
        RECT 107.575 47.565 108.075 47.735 ;
        RECT 108.955 47.565 109.455 47.735 ;
        RECT 107.575 46.650 108.075 46.820 ;
        RECT 108.955 46.650 109.455 46.820 ;
        RECT 107.345 45.395 107.515 46.435 ;
        RECT 108.135 45.395 108.305 46.435 ;
        RECT 108.725 45.395 108.895 46.435 ;
        RECT 109.515 45.395 109.685 46.435 ;
        RECT 110.230 44.935 110.940 49.510 ;
        RECT 111.420 44.940 112.130 49.515 ;
        RECT 112.670 47.950 112.840 48.990 ;
        RECT 113.460 47.950 113.630 48.990 ;
        RECT 114.050 47.950 114.220 48.990 ;
        RECT 114.840 47.950 115.010 48.990 ;
        RECT 112.900 47.565 113.400 47.735 ;
        RECT 114.280 47.565 114.780 47.735 ;
        RECT 112.900 46.650 113.400 46.820 ;
        RECT 114.280 46.650 114.780 46.820 ;
        RECT 112.670 45.395 112.840 46.435 ;
        RECT 113.460 45.395 113.630 46.435 ;
        RECT 114.050 45.395 114.220 46.435 ;
        RECT 114.840 45.395 115.010 46.435 ;
        RECT 115.555 44.935 116.265 49.510 ;
        RECT 116.755 44.940 117.465 49.515 ;
        RECT 118.005 47.950 118.175 48.990 ;
        RECT 118.795 47.950 118.965 48.990 ;
        RECT 119.385 47.950 119.555 48.990 ;
        RECT 120.175 47.950 120.345 48.990 ;
        RECT 118.235 47.565 118.735 47.735 ;
        RECT 119.615 47.565 120.115 47.735 ;
        RECT 118.235 46.650 118.735 46.820 ;
        RECT 119.615 46.650 120.115 46.820 ;
        RECT 118.005 45.395 118.175 46.435 ;
        RECT 118.795 45.395 118.965 46.435 ;
        RECT 119.385 45.395 119.555 46.435 ;
        RECT 120.175 45.395 120.345 46.435 ;
        RECT 120.890 44.935 121.600 49.510 ;
        RECT 122.080 44.955 122.790 49.530 ;
        RECT 123.330 47.950 123.500 48.990 ;
        RECT 124.120 47.950 124.290 48.990 ;
        RECT 124.710 47.950 124.880 48.990 ;
        RECT 125.500 47.950 125.670 48.990 ;
        RECT 123.330 45.395 123.500 46.435 ;
        RECT 124.120 45.395 124.290 46.435 ;
        RECT 124.710 45.395 124.880 46.435 ;
        RECT 125.500 45.395 125.670 46.435 ;
        RECT 126.215 44.955 126.925 49.530 ;
        RECT 14.565 44.485 20.400 44.655 ;
        RECT 16.175 44.470 20.400 44.485 ;
        RECT 14.645 44.265 15.945 44.295 ;
        RECT 12.130 44.060 12.685 44.230 ;
        RECT 12.455 43.820 12.685 44.060 ;
        RECT 13.600 44.030 20.050 44.265 ;
        RECT 12.090 42.990 12.685 43.820 ;
        RECT 14.485 43.845 19.515 43.850 ;
        RECT 20.230 43.845 20.400 44.470 ;
        RECT 32.725 43.950 32.895 44.640 ;
        RECT 33.515 43.950 33.685 44.640 ;
        RECT 34.105 43.950 34.275 44.640 ;
        RECT 34.895 43.950 35.065 44.640 ;
        RECT 38.050 43.950 38.220 44.640 ;
        RECT 38.840 43.950 39.010 44.640 ;
        RECT 39.430 43.950 39.600 44.640 ;
        RECT 40.220 43.950 40.390 44.640 ;
        RECT 43.385 43.950 43.555 44.640 ;
        RECT 44.175 43.950 44.345 44.640 ;
        RECT 44.765 43.950 44.935 44.640 ;
        RECT 45.555 43.950 45.725 44.640 ;
        RECT 48.710 43.950 48.880 44.640 ;
        RECT 49.500 43.950 49.670 44.640 ;
        RECT 50.090 43.950 50.260 44.640 ;
        RECT 50.880 43.950 51.050 44.640 ;
        RECT 54.045 43.950 54.215 44.640 ;
        RECT 54.835 43.950 55.005 44.640 ;
        RECT 55.425 43.950 55.595 44.640 ;
        RECT 56.215 43.950 56.385 44.640 ;
        RECT 59.370 43.950 59.540 44.640 ;
        RECT 60.160 43.950 60.330 44.640 ;
        RECT 60.750 43.950 60.920 44.640 ;
        RECT 61.540 43.950 61.710 44.640 ;
        RECT 64.705 43.950 64.875 44.640 ;
        RECT 65.495 43.950 65.665 44.640 ;
        RECT 66.085 43.950 66.255 44.640 ;
        RECT 66.875 43.950 67.045 44.640 ;
        RECT 70.030 43.950 70.200 44.640 ;
        RECT 70.820 43.950 70.990 44.640 ;
        RECT 71.410 43.950 71.580 44.640 ;
        RECT 72.200 43.950 72.370 44.640 ;
        RECT 75.365 43.950 75.535 44.640 ;
        RECT 76.155 43.950 76.325 44.640 ;
        RECT 76.745 43.950 76.915 44.640 ;
        RECT 77.535 43.950 77.705 44.640 ;
        RECT 80.690 43.950 80.860 44.640 ;
        RECT 81.480 43.950 81.650 44.640 ;
        RECT 82.070 43.950 82.240 44.640 ;
        RECT 82.860 43.950 83.030 44.640 ;
        RECT 86.025 43.950 86.195 44.640 ;
        RECT 86.815 43.950 86.985 44.640 ;
        RECT 87.405 43.950 87.575 44.640 ;
        RECT 88.195 43.950 88.365 44.640 ;
        RECT 91.350 43.950 91.520 44.640 ;
        RECT 92.140 43.950 92.310 44.640 ;
        RECT 92.730 43.950 92.900 44.640 ;
        RECT 93.520 43.950 93.690 44.640 ;
        RECT 96.685 43.950 96.855 44.640 ;
        RECT 97.475 43.950 97.645 44.640 ;
        RECT 98.065 43.950 98.235 44.640 ;
        RECT 98.855 43.950 99.025 44.640 ;
        RECT 102.010 43.950 102.180 44.640 ;
        RECT 102.800 43.950 102.970 44.640 ;
        RECT 103.390 43.950 103.560 44.640 ;
        RECT 104.180 43.950 104.350 44.640 ;
        RECT 107.345 43.950 107.515 44.640 ;
        RECT 108.135 43.950 108.305 44.640 ;
        RECT 108.725 43.950 108.895 44.640 ;
        RECT 109.515 43.950 109.685 44.640 ;
        RECT 112.670 43.950 112.840 44.640 ;
        RECT 113.460 43.950 113.630 44.640 ;
        RECT 114.050 43.950 114.220 44.640 ;
        RECT 114.840 43.950 115.010 44.640 ;
        RECT 118.005 43.950 118.175 44.640 ;
        RECT 118.795 43.950 118.965 44.640 ;
        RECT 119.385 43.950 119.555 44.640 ;
        RECT 120.175 43.950 120.345 44.640 ;
        RECT 123.330 43.950 123.500 44.640 ;
        RECT 124.120 43.950 124.290 44.640 ;
        RECT 124.710 43.950 124.880 44.640 ;
        RECT 125.500 43.950 125.670 44.640 ;
        RECT 14.485 43.680 20.400 43.845 ;
        RECT 14.485 43.180 14.695 43.680 ;
        RECT 16.045 43.675 20.400 43.680 ;
        RECT 16.045 43.665 20.260 43.675 ;
        RECT 16.045 43.180 16.255 43.665 ;
        RECT 17.605 43.180 17.815 43.665 ;
        RECT 19.205 43.180 19.855 43.665 ;
        RECT 38.280 43.610 38.780 43.780 ;
        RECT 39.660 43.610 40.160 43.780 ;
        RECT 43.615 43.610 44.115 43.780 ;
        RECT 44.995 43.610 45.495 43.780 ;
        RECT 48.940 43.610 49.440 43.780 ;
        RECT 50.320 43.610 50.820 43.780 ;
        RECT 54.275 43.610 54.775 43.780 ;
        RECT 55.655 43.610 56.155 43.780 ;
        RECT 59.600 43.610 60.100 43.780 ;
        RECT 60.980 43.610 61.480 43.780 ;
        RECT 64.935 43.610 65.435 43.780 ;
        RECT 66.315 43.610 66.815 43.780 ;
        RECT 70.260 43.610 70.760 43.780 ;
        RECT 71.640 43.610 72.140 43.780 ;
        RECT 75.595 43.610 76.095 43.780 ;
        RECT 76.975 43.610 77.475 43.780 ;
        RECT 80.920 43.610 81.420 43.780 ;
        RECT 82.300 43.610 82.800 43.780 ;
        RECT 86.255 43.610 86.755 43.780 ;
        RECT 87.635 43.610 88.135 43.780 ;
        RECT 91.580 43.610 92.080 43.780 ;
        RECT 92.960 43.610 93.460 43.780 ;
        RECT 96.915 43.610 97.415 43.780 ;
        RECT 98.295 43.610 98.795 43.780 ;
        RECT 102.240 43.610 102.740 43.780 ;
        RECT 103.620 43.610 104.120 43.780 ;
        RECT 107.575 43.610 108.075 43.780 ;
        RECT 108.955 43.610 109.455 43.780 ;
        RECT 112.900 43.610 113.400 43.780 ;
        RECT 114.280 43.610 114.780 43.780 ;
        RECT 118.235 43.610 118.735 43.780 ;
        RECT 119.615 43.610 120.115 43.780 ;
        RECT 38.280 43.070 38.780 43.240 ;
        RECT 39.660 43.070 40.160 43.240 ;
        RECT 43.615 43.070 44.115 43.240 ;
        RECT 44.995 43.070 45.495 43.240 ;
        RECT 48.940 43.070 49.440 43.240 ;
        RECT 50.320 43.070 50.820 43.240 ;
        RECT 54.275 43.070 54.775 43.240 ;
        RECT 55.655 43.070 56.155 43.240 ;
        RECT 59.600 43.070 60.100 43.240 ;
        RECT 60.980 43.070 61.480 43.240 ;
        RECT 64.935 43.070 65.435 43.240 ;
        RECT 66.315 43.070 66.815 43.240 ;
        RECT 70.260 43.070 70.760 43.240 ;
        RECT 71.640 43.070 72.140 43.240 ;
        RECT 75.595 43.070 76.095 43.240 ;
        RECT 76.975 43.070 77.475 43.240 ;
        RECT 80.920 43.070 81.420 43.240 ;
        RECT 82.300 43.070 82.800 43.240 ;
        RECT 86.255 43.070 86.755 43.240 ;
        RECT 87.635 43.070 88.135 43.240 ;
        RECT 91.580 43.070 92.080 43.240 ;
        RECT 92.960 43.070 93.460 43.240 ;
        RECT 96.915 43.070 97.415 43.240 ;
        RECT 98.295 43.070 98.795 43.240 ;
        RECT 102.240 43.070 102.740 43.240 ;
        RECT 103.620 43.070 104.120 43.240 ;
        RECT 107.575 43.070 108.075 43.240 ;
        RECT 108.955 43.070 109.455 43.240 ;
        RECT 112.900 43.070 113.400 43.240 ;
        RECT 114.280 43.070 114.780 43.240 ;
        RECT 118.235 43.070 118.735 43.240 ;
        RECT 119.615 43.070 120.115 43.240 ;
        RECT 32.725 42.210 32.895 42.900 ;
        RECT 33.515 42.210 33.685 42.900 ;
        RECT 34.105 42.210 34.275 42.900 ;
        RECT 34.895 42.210 35.065 42.900 ;
        RECT 38.050 42.210 38.220 42.900 ;
        RECT 38.840 42.210 39.010 42.900 ;
        RECT 39.430 42.210 39.600 42.900 ;
        RECT 40.220 42.210 40.390 42.900 ;
        RECT 43.385 42.210 43.555 42.900 ;
        RECT 44.175 42.210 44.345 42.900 ;
        RECT 44.765 42.210 44.935 42.900 ;
        RECT 45.555 42.210 45.725 42.900 ;
        RECT 48.710 42.210 48.880 42.900 ;
        RECT 49.500 42.210 49.670 42.900 ;
        RECT 50.090 42.210 50.260 42.900 ;
        RECT 50.880 42.210 51.050 42.900 ;
        RECT 54.045 42.210 54.215 42.900 ;
        RECT 54.835 42.210 55.005 42.900 ;
        RECT 55.425 42.210 55.595 42.900 ;
        RECT 56.215 42.210 56.385 42.900 ;
        RECT 59.370 42.210 59.540 42.900 ;
        RECT 60.160 42.210 60.330 42.900 ;
        RECT 60.750 42.210 60.920 42.900 ;
        RECT 61.540 42.210 61.710 42.900 ;
        RECT 64.705 42.210 64.875 42.900 ;
        RECT 65.495 42.210 65.665 42.900 ;
        RECT 66.085 42.210 66.255 42.900 ;
        RECT 66.875 42.210 67.045 42.900 ;
        RECT 70.030 42.210 70.200 42.900 ;
        RECT 70.820 42.210 70.990 42.900 ;
        RECT 71.410 42.210 71.580 42.900 ;
        RECT 72.200 42.210 72.370 42.900 ;
        RECT 75.365 42.210 75.535 42.900 ;
        RECT 76.155 42.210 76.325 42.900 ;
        RECT 76.745 42.210 76.915 42.900 ;
        RECT 77.535 42.210 77.705 42.900 ;
        RECT 80.690 42.210 80.860 42.900 ;
        RECT 81.480 42.210 81.650 42.900 ;
        RECT 82.070 42.210 82.240 42.900 ;
        RECT 82.860 42.210 83.030 42.900 ;
        RECT 86.025 42.210 86.195 42.900 ;
        RECT 86.815 42.210 86.985 42.900 ;
        RECT 87.405 42.210 87.575 42.900 ;
        RECT 88.195 42.210 88.365 42.900 ;
        RECT 91.350 42.210 91.520 42.900 ;
        RECT 92.140 42.210 92.310 42.900 ;
        RECT 92.730 42.210 92.900 42.900 ;
        RECT 93.520 42.210 93.690 42.900 ;
        RECT 96.685 42.210 96.855 42.900 ;
        RECT 97.475 42.210 97.645 42.900 ;
        RECT 98.065 42.210 98.235 42.900 ;
        RECT 98.855 42.210 99.025 42.900 ;
        RECT 102.010 42.210 102.180 42.900 ;
        RECT 102.800 42.210 102.970 42.900 ;
        RECT 103.390 42.210 103.560 42.900 ;
        RECT 104.180 42.210 104.350 42.900 ;
        RECT 107.345 42.210 107.515 42.900 ;
        RECT 108.135 42.210 108.305 42.900 ;
        RECT 108.725 42.210 108.895 42.900 ;
        RECT 109.515 42.210 109.685 42.900 ;
        RECT 112.670 42.210 112.840 42.900 ;
        RECT 113.460 42.210 113.630 42.900 ;
        RECT 114.050 42.210 114.220 42.900 ;
        RECT 114.840 42.210 115.010 42.900 ;
        RECT 118.005 42.210 118.175 42.900 ;
        RECT 118.795 42.210 118.965 42.900 ;
        RECT 119.385 42.210 119.555 42.900 ;
        RECT 120.175 42.210 120.345 42.900 ;
        RECT 123.330 42.210 123.500 42.900 ;
        RECT 124.120 42.210 124.290 42.900 ;
        RECT 124.710 42.210 124.880 42.900 ;
        RECT 125.500 42.210 125.670 42.900 ;
        RECT 2.825 40.305 3.155 41.855 ;
        RECT 4.385 40.305 4.715 41.855 ;
        RECT 5.945 40.305 6.275 41.935 ;
        RECT 8.845 40.865 9.175 41.935 ;
        RECT 10.450 41.035 10.780 41.935 ;
        RECT 11.930 41.220 12.180 41.955 ;
        RECT 13.490 41.220 14.075 41.955 ;
        RECT 11.930 41.050 14.075 41.220 ;
        RECT 15.925 41.225 16.135 41.720 ;
        RECT 17.485 41.225 17.695 41.720 ;
        RECT 19.045 41.225 19.255 41.720 ;
        RECT 20.645 41.225 21.295 41.720 ;
        RECT 15.925 41.050 21.840 41.225 ;
        RECT 7.990 40.305 8.320 40.865 ;
        RECT 2.825 39.975 8.320 40.305 ;
        RECT 3.215 37.365 3.505 39.805 ;
        RECT 6.515 37.775 6.845 39.975 ;
        RECT 7.990 39.515 8.320 39.975 ;
        RECT 8.845 40.535 10.370 40.865 ;
        RECT 7.015 38.780 7.825 39.110 ;
        RECT 7.495 38.115 7.825 38.780 ;
        RECT 8.845 38.715 9.175 40.535 ;
        RECT 10.540 40.365 10.780 41.035 ;
        RECT 13.905 40.900 14.075 41.050 ;
        RECT 13.905 40.870 14.605 40.900 ;
        RECT 11.015 40.700 13.725 40.870 ;
        RECT 13.905 40.635 21.490 40.870 ;
        RECT 13.905 40.520 15.710 40.635 ;
        RECT 10.450 38.715 10.780 40.365 ;
        RECT 11.930 40.350 15.710 40.520 ;
        RECT 21.670 40.420 21.840 41.050 ;
        RECT 16.045 40.415 21.840 40.420 ;
        RECT 11.930 38.695 12.260 40.350 ;
        RECT 13.570 38.695 13.820 40.350 ;
        RECT 16.005 40.245 21.840 40.415 ;
        RECT 16.005 39.005 16.335 40.245 ;
        RECT 17.565 39.005 17.895 40.245 ;
        RECT 19.125 39.005 19.455 40.245 ;
        RECT 20.685 39.005 21.015 40.245 ;
        RECT 6.515 37.445 7.325 37.775 ;
        RECT 3.215 37.075 3.595 37.365 ;
        RECT 3.305 36.305 3.595 37.075 ;
        RECT 4.205 36.785 4.515 37.215 ;
        RECT 6.995 37.105 7.325 37.445 ;
        RECT 7.495 37.705 8.165 38.115 ;
        RECT 7.495 36.785 7.825 37.705 ;
        RECT 4.205 36.475 6.120 36.785 ;
        RECT 4.810 36.455 6.120 36.475 ;
        RECT 6.290 36.455 9.740 36.785 ;
        RECT 3.305 36.055 4.640 36.305 ;
        RECT 3.305 35.045 3.595 36.055 ;
        RECT 4.810 35.885 5.140 36.455 ;
        RECT 4.205 35.555 5.140 35.885 ;
        RECT 4.205 35.045 4.515 35.555 ;
        RECT 6.290 34.905 6.620 36.455 ;
        RECT 7.850 34.905 8.180 36.455 ;
        RECT 9.410 34.825 9.740 36.455 ;
        RECT 11.015 35.860 11.960 36.190 ;
        RECT 12.130 36.090 12.380 38.065 ;
        RECT 14.565 36.515 14.895 37.755 ;
        RECT 16.125 36.515 16.455 37.755 ;
        RECT 17.685 36.515 18.015 37.755 ;
        RECT 19.245 36.515 19.575 37.755 ;
        RECT 31.475 37.420 32.185 41.995 ;
        RECT 32.725 40.415 32.895 41.455 ;
        RECT 33.515 40.415 33.685 41.455 ;
        RECT 34.105 40.415 34.275 41.455 ;
        RECT 34.895 40.415 35.065 41.455 ;
        RECT 32.725 37.860 32.895 38.900 ;
        RECT 33.515 37.860 33.685 38.900 ;
        RECT 34.105 37.860 34.275 38.900 ;
        RECT 34.895 37.860 35.065 38.900 ;
        RECT 35.610 37.420 36.320 41.995 ;
        RECT 36.800 37.405 37.510 41.980 ;
        RECT 38.050 40.415 38.220 41.455 ;
        RECT 38.840 40.415 39.010 41.455 ;
        RECT 39.430 40.415 39.600 41.455 ;
        RECT 40.220 40.415 40.390 41.455 ;
        RECT 38.280 40.030 38.780 40.200 ;
        RECT 39.660 40.030 40.160 40.200 ;
        RECT 38.280 39.115 38.780 39.285 ;
        RECT 39.660 39.115 40.160 39.285 ;
        RECT 38.050 37.860 38.220 38.900 ;
        RECT 38.840 37.860 39.010 38.900 ;
        RECT 39.430 37.860 39.600 38.900 ;
        RECT 40.220 37.860 40.390 38.900 ;
        RECT 40.935 37.400 41.645 41.975 ;
        RECT 42.135 37.405 42.845 41.980 ;
        RECT 43.385 40.415 43.555 41.455 ;
        RECT 44.175 40.415 44.345 41.455 ;
        RECT 44.765 40.415 44.935 41.455 ;
        RECT 45.555 40.415 45.725 41.455 ;
        RECT 43.615 40.030 44.115 40.200 ;
        RECT 44.995 40.030 45.495 40.200 ;
        RECT 43.615 39.115 44.115 39.285 ;
        RECT 44.995 39.115 45.495 39.285 ;
        RECT 43.385 37.860 43.555 38.900 ;
        RECT 44.175 37.860 44.345 38.900 ;
        RECT 44.765 37.860 44.935 38.900 ;
        RECT 45.555 37.860 45.725 38.900 ;
        RECT 46.270 37.400 46.980 41.975 ;
        RECT 47.460 37.405 48.170 41.980 ;
        RECT 48.710 40.415 48.880 41.455 ;
        RECT 49.500 40.415 49.670 41.455 ;
        RECT 50.090 40.415 50.260 41.455 ;
        RECT 50.880 40.415 51.050 41.455 ;
        RECT 48.940 40.030 49.440 40.200 ;
        RECT 50.320 40.030 50.820 40.200 ;
        RECT 48.940 39.115 49.440 39.285 ;
        RECT 50.320 39.115 50.820 39.285 ;
        RECT 48.710 37.860 48.880 38.900 ;
        RECT 49.500 37.860 49.670 38.900 ;
        RECT 50.090 37.860 50.260 38.900 ;
        RECT 50.880 37.860 51.050 38.900 ;
        RECT 51.595 37.400 52.305 41.975 ;
        RECT 52.795 37.405 53.505 41.980 ;
        RECT 54.045 40.415 54.215 41.455 ;
        RECT 54.835 40.415 55.005 41.455 ;
        RECT 55.425 40.415 55.595 41.455 ;
        RECT 56.215 40.415 56.385 41.455 ;
        RECT 54.275 40.030 54.775 40.200 ;
        RECT 55.655 40.030 56.155 40.200 ;
        RECT 54.275 39.115 54.775 39.285 ;
        RECT 55.655 39.115 56.155 39.285 ;
        RECT 54.045 37.860 54.215 38.900 ;
        RECT 54.835 37.860 55.005 38.900 ;
        RECT 55.425 37.860 55.595 38.900 ;
        RECT 56.215 37.860 56.385 38.900 ;
        RECT 56.930 37.400 57.640 41.975 ;
        RECT 58.120 37.405 58.830 41.980 ;
        RECT 59.370 40.415 59.540 41.455 ;
        RECT 60.160 40.415 60.330 41.455 ;
        RECT 60.750 40.415 60.920 41.455 ;
        RECT 61.540 40.415 61.710 41.455 ;
        RECT 59.600 40.030 60.100 40.200 ;
        RECT 60.980 40.030 61.480 40.200 ;
        RECT 59.600 39.115 60.100 39.285 ;
        RECT 60.980 39.115 61.480 39.285 ;
        RECT 59.370 37.860 59.540 38.900 ;
        RECT 60.160 37.860 60.330 38.900 ;
        RECT 60.750 37.860 60.920 38.900 ;
        RECT 61.540 37.860 61.710 38.900 ;
        RECT 62.255 37.400 62.965 41.975 ;
        RECT 63.455 37.405 64.165 41.980 ;
        RECT 64.705 40.415 64.875 41.455 ;
        RECT 65.495 40.415 65.665 41.455 ;
        RECT 66.085 40.415 66.255 41.455 ;
        RECT 66.875 40.415 67.045 41.455 ;
        RECT 64.935 40.030 65.435 40.200 ;
        RECT 66.315 40.030 66.815 40.200 ;
        RECT 64.935 39.115 65.435 39.285 ;
        RECT 66.315 39.115 66.815 39.285 ;
        RECT 64.705 37.860 64.875 38.900 ;
        RECT 65.495 37.860 65.665 38.900 ;
        RECT 66.085 37.860 66.255 38.900 ;
        RECT 66.875 37.860 67.045 38.900 ;
        RECT 67.590 37.400 68.300 41.975 ;
        RECT 68.780 37.405 69.490 41.980 ;
        RECT 70.030 40.415 70.200 41.455 ;
        RECT 70.820 40.415 70.990 41.455 ;
        RECT 71.410 40.415 71.580 41.455 ;
        RECT 72.200 40.415 72.370 41.455 ;
        RECT 70.260 40.030 70.760 40.200 ;
        RECT 71.640 40.030 72.140 40.200 ;
        RECT 70.260 39.115 70.760 39.285 ;
        RECT 71.640 39.115 72.140 39.285 ;
        RECT 70.030 37.860 70.200 38.900 ;
        RECT 70.820 37.860 70.990 38.900 ;
        RECT 71.410 37.860 71.580 38.900 ;
        RECT 72.200 37.860 72.370 38.900 ;
        RECT 72.915 37.400 73.625 41.975 ;
        RECT 74.115 37.405 74.825 41.980 ;
        RECT 75.365 40.415 75.535 41.455 ;
        RECT 76.155 40.415 76.325 41.455 ;
        RECT 76.745 40.415 76.915 41.455 ;
        RECT 77.535 40.415 77.705 41.455 ;
        RECT 75.595 40.030 76.095 40.200 ;
        RECT 76.975 40.030 77.475 40.200 ;
        RECT 75.595 39.115 76.095 39.285 ;
        RECT 76.975 39.115 77.475 39.285 ;
        RECT 75.365 37.860 75.535 38.900 ;
        RECT 76.155 37.860 76.325 38.900 ;
        RECT 76.745 37.860 76.915 38.900 ;
        RECT 77.535 37.860 77.705 38.900 ;
        RECT 78.250 37.400 78.960 41.975 ;
        RECT 79.440 37.405 80.150 41.980 ;
        RECT 80.690 40.415 80.860 41.455 ;
        RECT 81.480 40.415 81.650 41.455 ;
        RECT 82.070 40.415 82.240 41.455 ;
        RECT 82.860 40.415 83.030 41.455 ;
        RECT 80.920 40.030 81.420 40.200 ;
        RECT 82.300 40.030 82.800 40.200 ;
        RECT 80.920 39.115 81.420 39.285 ;
        RECT 82.300 39.115 82.800 39.285 ;
        RECT 80.690 37.860 80.860 38.900 ;
        RECT 81.480 37.860 81.650 38.900 ;
        RECT 82.070 37.860 82.240 38.900 ;
        RECT 82.860 37.860 83.030 38.900 ;
        RECT 83.575 37.400 84.285 41.975 ;
        RECT 84.775 37.405 85.485 41.980 ;
        RECT 86.025 40.415 86.195 41.455 ;
        RECT 86.815 40.415 86.985 41.455 ;
        RECT 87.405 40.415 87.575 41.455 ;
        RECT 88.195 40.415 88.365 41.455 ;
        RECT 86.255 40.030 86.755 40.200 ;
        RECT 87.635 40.030 88.135 40.200 ;
        RECT 86.255 39.115 86.755 39.285 ;
        RECT 87.635 39.115 88.135 39.285 ;
        RECT 86.025 37.860 86.195 38.900 ;
        RECT 86.815 37.860 86.985 38.900 ;
        RECT 87.405 37.860 87.575 38.900 ;
        RECT 88.195 37.860 88.365 38.900 ;
        RECT 88.910 37.400 89.620 41.975 ;
        RECT 90.100 37.405 90.810 41.980 ;
        RECT 91.350 40.415 91.520 41.455 ;
        RECT 92.140 40.415 92.310 41.455 ;
        RECT 92.730 40.415 92.900 41.455 ;
        RECT 93.520 40.415 93.690 41.455 ;
        RECT 91.580 40.030 92.080 40.200 ;
        RECT 92.960 40.030 93.460 40.200 ;
        RECT 91.580 39.115 92.080 39.285 ;
        RECT 92.960 39.115 93.460 39.285 ;
        RECT 91.350 37.860 91.520 38.900 ;
        RECT 92.140 37.860 92.310 38.900 ;
        RECT 92.730 37.860 92.900 38.900 ;
        RECT 93.520 37.860 93.690 38.900 ;
        RECT 94.235 37.400 94.945 41.975 ;
        RECT 95.435 37.405 96.145 41.980 ;
        RECT 96.685 40.415 96.855 41.455 ;
        RECT 97.475 40.415 97.645 41.455 ;
        RECT 98.065 40.415 98.235 41.455 ;
        RECT 98.855 40.415 99.025 41.455 ;
        RECT 96.915 40.030 97.415 40.200 ;
        RECT 98.295 40.030 98.795 40.200 ;
        RECT 96.915 39.115 97.415 39.285 ;
        RECT 98.295 39.115 98.795 39.285 ;
        RECT 96.685 37.860 96.855 38.900 ;
        RECT 97.475 37.860 97.645 38.900 ;
        RECT 98.065 37.860 98.235 38.900 ;
        RECT 98.855 37.860 99.025 38.900 ;
        RECT 99.570 37.400 100.280 41.975 ;
        RECT 100.760 37.405 101.470 41.980 ;
        RECT 102.010 40.415 102.180 41.455 ;
        RECT 102.800 40.415 102.970 41.455 ;
        RECT 103.390 40.415 103.560 41.455 ;
        RECT 104.180 40.415 104.350 41.455 ;
        RECT 102.240 40.030 102.740 40.200 ;
        RECT 103.620 40.030 104.120 40.200 ;
        RECT 102.240 39.115 102.740 39.285 ;
        RECT 103.620 39.115 104.120 39.285 ;
        RECT 102.010 37.860 102.180 38.900 ;
        RECT 102.800 37.860 102.970 38.900 ;
        RECT 103.390 37.860 103.560 38.900 ;
        RECT 104.180 37.860 104.350 38.900 ;
        RECT 104.895 37.400 105.605 41.975 ;
        RECT 106.095 37.405 106.805 41.980 ;
        RECT 107.345 40.415 107.515 41.455 ;
        RECT 108.135 40.415 108.305 41.455 ;
        RECT 108.725 40.415 108.895 41.455 ;
        RECT 109.515 40.415 109.685 41.455 ;
        RECT 107.575 40.030 108.075 40.200 ;
        RECT 108.955 40.030 109.455 40.200 ;
        RECT 107.575 39.115 108.075 39.285 ;
        RECT 108.955 39.115 109.455 39.285 ;
        RECT 107.345 37.860 107.515 38.900 ;
        RECT 108.135 37.860 108.305 38.900 ;
        RECT 108.725 37.860 108.895 38.900 ;
        RECT 109.515 37.860 109.685 38.900 ;
        RECT 110.230 37.400 110.940 41.975 ;
        RECT 111.420 37.405 112.130 41.980 ;
        RECT 112.670 40.415 112.840 41.455 ;
        RECT 113.460 40.415 113.630 41.455 ;
        RECT 114.050 40.415 114.220 41.455 ;
        RECT 114.840 40.415 115.010 41.455 ;
        RECT 112.900 40.030 113.400 40.200 ;
        RECT 114.280 40.030 114.780 40.200 ;
        RECT 112.900 39.115 113.400 39.285 ;
        RECT 114.280 39.115 114.780 39.285 ;
        RECT 112.670 37.860 112.840 38.900 ;
        RECT 113.460 37.860 113.630 38.900 ;
        RECT 114.050 37.860 114.220 38.900 ;
        RECT 114.840 37.860 115.010 38.900 ;
        RECT 115.555 37.400 116.265 41.975 ;
        RECT 116.755 37.405 117.465 41.980 ;
        RECT 118.005 40.415 118.175 41.455 ;
        RECT 118.795 40.415 118.965 41.455 ;
        RECT 119.385 40.415 119.555 41.455 ;
        RECT 120.175 40.415 120.345 41.455 ;
        RECT 118.235 40.030 118.735 40.200 ;
        RECT 119.615 40.030 120.115 40.200 ;
        RECT 118.235 39.115 118.735 39.285 ;
        RECT 119.615 39.115 120.115 39.285 ;
        RECT 118.005 37.860 118.175 38.900 ;
        RECT 118.795 37.860 118.965 38.900 ;
        RECT 119.385 37.860 119.555 38.900 ;
        RECT 120.175 37.860 120.345 38.900 ;
        RECT 120.890 37.400 121.600 41.975 ;
        RECT 122.080 37.420 122.790 41.995 ;
        RECT 123.330 40.415 123.500 41.455 ;
        RECT 124.120 40.415 124.290 41.455 ;
        RECT 124.710 40.415 124.880 41.455 ;
        RECT 125.500 40.415 125.670 41.455 ;
        RECT 123.330 37.860 123.500 38.900 ;
        RECT 124.120 37.860 124.290 38.900 ;
        RECT 124.710 37.860 124.880 38.900 ;
        RECT 125.500 37.860 125.670 38.900 ;
        RECT 126.215 37.420 126.925 41.995 ;
        RECT 14.565 36.345 20.400 36.515 ;
        RECT 32.725 36.415 32.895 37.105 ;
        RECT 33.515 36.415 33.685 37.105 ;
        RECT 34.105 36.415 34.275 37.105 ;
        RECT 34.895 36.415 35.065 37.105 ;
        RECT 38.050 36.415 38.220 37.105 ;
        RECT 38.840 36.415 39.010 37.105 ;
        RECT 39.430 36.415 39.600 37.105 ;
        RECT 40.220 36.415 40.390 37.105 ;
        RECT 43.385 36.415 43.555 37.105 ;
        RECT 44.175 36.415 44.345 37.105 ;
        RECT 44.765 36.415 44.935 37.105 ;
        RECT 45.555 36.415 45.725 37.105 ;
        RECT 48.710 36.415 48.880 37.105 ;
        RECT 49.500 36.415 49.670 37.105 ;
        RECT 50.090 36.415 50.260 37.105 ;
        RECT 50.880 36.415 51.050 37.105 ;
        RECT 54.045 36.415 54.215 37.105 ;
        RECT 54.835 36.415 55.005 37.105 ;
        RECT 55.425 36.415 55.595 37.105 ;
        RECT 56.215 36.415 56.385 37.105 ;
        RECT 59.370 36.415 59.540 37.105 ;
        RECT 60.160 36.415 60.330 37.105 ;
        RECT 60.750 36.415 60.920 37.105 ;
        RECT 61.540 36.415 61.710 37.105 ;
        RECT 64.705 36.415 64.875 37.105 ;
        RECT 65.495 36.415 65.665 37.105 ;
        RECT 66.085 36.415 66.255 37.105 ;
        RECT 66.875 36.415 67.045 37.105 ;
        RECT 70.030 36.415 70.200 37.105 ;
        RECT 70.820 36.415 70.990 37.105 ;
        RECT 71.410 36.415 71.580 37.105 ;
        RECT 72.200 36.415 72.370 37.105 ;
        RECT 75.365 36.415 75.535 37.105 ;
        RECT 76.155 36.415 76.325 37.105 ;
        RECT 76.745 36.415 76.915 37.105 ;
        RECT 77.535 36.415 77.705 37.105 ;
        RECT 80.690 36.415 80.860 37.105 ;
        RECT 81.480 36.415 81.650 37.105 ;
        RECT 82.070 36.415 82.240 37.105 ;
        RECT 82.860 36.415 83.030 37.105 ;
        RECT 86.025 36.415 86.195 37.105 ;
        RECT 86.815 36.415 86.985 37.105 ;
        RECT 87.405 36.415 87.575 37.105 ;
        RECT 88.195 36.415 88.365 37.105 ;
        RECT 91.350 36.415 91.520 37.105 ;
        RECT 92.140 36.415 92.310 37.105 ;
        RECT 92.730 36.415 92.900 37.105 ;
        RECT 93.520 36.415 93.690 37.105 ;
        RECT 96.685 36.415 96.855 37.105 ;
        RECT 97.475 36.415 97.645 37.105 ;
        RECT 98.065 36.415 98.235 37.105 ;
        RECT 98.855 36.415 99.025 37.105 ;
        RECT 102.010 36.415 102.180 37.105 ;
        RECT 102.800 36.415 102.970 37.105 ;
        RECT 103.390 36.415 103.560 37.105 ;
        RECT 104.180 36.415 104.350 37.105 ;
        RECT 107.345 36.415 107.515 37.105 ;
        RECT 108.135 36.415 108.305 37.105 ;
        RECT 108.725 36.415 108.895 37.105 ;
        RECT 109.515 36.415 109.685 37.105 ;
        RECT 112.670 36.415 112.840 37.105 ;
        RECT 113.460 36.415 113.630 37.105 ;
        RECT 114.050 36.415 114.220 37.105 ;
        RECT 114.840 36.415 115.010 37.105 ;
        RECT 118.005 36.415 118.175 37.105 ;
        RECT 118.795 36.415 118.965 37.105 ;
        RECT 119.385 36.415 119.555 37.105 ;
        RECT 120.175 36.415 120.345 37.105 ;
        RECT 123.330 36.415 123.500 37.105 ;
        RECT 124.120 36.415 124.290 37.105 ;
        RECT 124.710 36.415 124.880 37.105 ;
        RECT 125.500 36.415 125.670 37.105 ;
        RECT 16.175 36.330 20.400 36.345 ;
        RECT 14.645 36.125 15.945 36.155 ;
        RECT 12.130 35.920 12.685 36.090 ;
        RECT 12.455 35.680 12.685 35.920 ;
        RECT 13.600 35.890 20.050 36.125 ;
        RECT 12.090 34.850 12.685 35.680 ;
        RECT 14.485 35.705 19.515 35.710 ;
        RECT 20.230 35.705 20.400 36.330 ;
        RECT 38.280 36.075 38.780 36.245 ;
        RECT 39.660 36.075 40.160 36.245 ;
        RECT 43.615 36.075 44.115 36.245 ;
        RECT 44.995 36.075 45.495 36.245 ;
        RECT 48.940 36.075 49.440 36.245 ;
        RECT 50.320 36.075 50.820 36.245 ;
        RECT 54.275 36.075 54.775 36.245 ;
        RECT 55.655 36.075 56.155 36.245 ;
        RECT 59.600 36.075 60.100 36.245 ;
        RECT 60.980 36.075 61.480 36.245 ;
        RECT 64.935 36.075 65.435 36.245 ;
        RECT 66.315 36.075 66.815 36.245 ;
        RECT 70.260 36.075 70.760 36.245 ;
        RECT 71.640 36.075 72.140 36.245 ;
        RECT 75.595 36.075 76.095 36.245 ;
        RECT 76.975 36.075 77.475 36.245 ;
        RECT 80.920 36.075 81.420 36.245 ;
        RECT 82.300 36.075 82.800 36.245 ;
        RECT 86.255 36.075 86.755 36.245 ;
        RECT 87.635 36.075 88.135 36.245 ;
        RECT 91.580 36.075 92.080 36.245 ;
        RECT 92.960 36.075 93.460 36.245 ;
        RECT 96.915 36.075 97.415 36.245 ;
        RECT 98.295 36.075 98.795 36.245 ;
        RECT 102.240 36.075 102.740 36.245 ;
        RECT 103.620 36.075 104.120 36.245 ;
        RECT 107.575 36.075 108.075 36.245 ;
        RECT 108.955 36.075 109.455 36.245 ;
        RECT 112.900 36.075 113.400 36.245 ;
        RECT 114.280 36.075 114.780 36.245 ;
        RECT 118.235 36.075 118.735 36.245 ;
        RECT 119.615 36.075 120.115 36.245 ;
        RECT 14.485 35.540 20.400 35.705 ;
        RECT 14.485 35.040 14.695 35.540 ;
        RECT 16.045 35.535 20.400 35.540 ;
        RECT 38.280 35.535 38.780 35.705 ;
        RECT 39.660 35.535 40.160 35.705 ;
        RECT 43.615 35.535 44.115 35.705 ;
        RECT 44.995 35.535 45.495 35.705 ;
        RECT 48.940 35.535 49.440 35.705 ;
        RECT 50.320 35.535 50.820 35.705 ;
        RECT 54.275 35.535 54.775 35.705 ;
        RECT 55.655 35.535 56.155 35.705 ;
        RECT 59.600 35.535 60.100 35.705 ;
        RECT 60.980 35.535 61.480 35.705 ;
        RECT 64.935 35.535 65.435 35.705 ;
        RECT 66.315 35.535 66.815 35.705 ;
        RECT 70.260 35.535 70.760 35.705 ;
        RECT 71.640 35.535 72.140 35.705 ;
        RECT 75.595 35.535 76.095 35.705 ;
        RECT 76.975 35.535 77.475 35.705 ;
        RECT 80.920 35.535 81.420 35.705 ;
        RECT 82.300 35.535 82.800 35.705 ;
        RECT 86.255 35.535 86.755 35.705 ;
        RECT 87.635 35.535 88.135 35.705 ;
        RECT 91.580 35.535 92.080 35.705 ;
        RECT 92.960 35.535 93.460 35.705 ;
        RECT 96.915 35.535 97.415 35.705 ;
        RECT 98.295 35.535 98.795 35.705 ;
        RECT 102.240 35.535 102.740 35.705 ;
        RECT 103.620 35.535 104.120 35.705 ;
        RECT 107.575 35.535 108.075 35.705 ;
        RECT 108.955 35.535 109.455 35.705 ;
        RECT 112.900 35.535 113.400 35.705 ;
        RECT 114.280 35.535 114.780 35.705 ;
        RECT 118.235 35.535 118.735 35.705 ;
        RECT 119.615 35.535 120.115 35.705 ;
        RECT 16.045 35.525 20.260 35.535 ;
        RECT 16.045 35.040 16.255 35.525 ;
        RECT 17.605 35.040 17.815 35.525 ;
        RECT 19.205 35.040 19.855 35.525 ;
        RECT 32.725 34.675 32.895 35.365 ;
        RECT 33.515 34.675 33.685 35.365 ;
        RECT 34.105 34.675 34.275 35.365 ;
        RECT 34.895 34.675 35.065 35.365 ;
        RECT 38.050 34.675 38.220 35.365 ;
        RECT 38.840 34.675 39.010 35.365 ;
        RECT 39.430 34.675 39.600 35.365 ;
        RECT 40.220 34.675 40.390 35.365 ;
        RECT 43.385 34.675 43.555 35.365 ;
        RECT 44.175 34.675 44.345 35.365 ;
        RECT 44.765 34.675 44.935 35.365 ;
        RECT 45.555 34.675 45.725 35.365 ;
        RECT 48.710 34.675 48.880 35.365 ;
        RECT 49.500 34.675 49.670 35.365 ;
        RECT 50.090 34.675 50.260 35.365 ;
        RECT 50.880 34.675 51.050 35.365 ;
        RECT 54.045 34.675 54.215 35.365 ;
        RECT 54.835 34.675 55.005 35.365 ;
        RECT 55.425 34.675 55.595 35.365 ;
        RECT 56.215 34.675 56.385 35.365 ;
        RECT 59.370 34.675 59.540 35.365 ;
        RECT 60.160 34.675 60.330 35.365 ;
        RECT 60.750 34.675 60.920 35.365 ;
        RECT 61.540 34.675 61.710 35.365 ;
        RECT 64.705 34.675 64.875 35.365 ;
        RECT 65.495 34.675 65.665 35.365 ;
        RECT 66.085 34.675 66.255 35.365 ;
        RECT 66.875 34.675 67.045 35.365 ;
        RECT 70.030 34.675 70.200 35.365 ;
        RECT 70.820 34.675 70.990 35.365 ;
        RECT 71.410 34.675 71.580 35.365 ;
        RECT 72.200 34.675 72.370 35.365 ;
        RECT 75.365 34.675 75.535 35.365 ;
        RECT 76.155 34.675 76.325 35.365 ;
        RECT 76.745 34.675 76.915 35.365 ;
        RECT 77.535 34.675 77.705 35.365 ;
        RECT 80.690 34.675 80.860 35.365 ;
        RECT 81.480 34.675 81.650 35.365 ;
        RECT 82.070 34.675 82.240 35.365 ;
        RECT 82.860 34.675 83.030 35.365 ;
        RECT 86.025 34.675 86.195 35.365 ;
        RECT 86.815 34.675 86.985 35.365 ;
        RECT 87.405 34.675 87.575 35.365 ;
        RECT 88.195 34.675 88.365 35.365 ;
        RECT 91.350 34.675 91.520 35.365 ;
        RECT 92.140 34.675 92.310 35.365 ;
        RECT 92.730 34.675 92.900 35.365 ;
        RECT 93.520 34.675 93.690 35.365 ;
        RECT 96.685 34.675 96.855 35.365 ;
        RECT 97.475 34.675 97.645 35.365 ;
        RECT 98.065 34.675 98.235 35.365 ;
        RECT 98.855 34.675 99.025 35.365 ;
        RECT 102.010 34.675 102.180 35.365 ;
        RECT 102.800 34.675 102.970 35.365 ;
        RECT 103.390 34.675 103.560 35.365 ;
        RECT 104.180 34.675 104.350 35.365 ;
        RECT 107.345 34.675 107.515 35.365 ;
        RECT 108.135 34.675 108.305 35.365 ;
        RECT 108.725 34.675 108.895 35.365 ;
        RECT 109.515 34.675 109.685 35.365 ;
        RECT 112.670 34.675 112.840 35.365 ;
        RECT 113.460 34.675 113.630 35.365 ;
        RECT 114.050 34.675 114.220 35.365 ;
        RECT 114.840 34.675 115.010 35.365 ;
        RECT 118.005 34.675 118.175 35.365 ;
        RECT 118.795 34.675 118.965 35.365 ;
        RECT 119.385 34.675 119.555 35.365 ;
        RECT 120.175 34.675 120.345 35.365 ;
        RECT 123.330 34.675 123.500 35.365 ;
        RECT 124.120 34.675 124.290 35.365 ;
        RECT 124.710 34.675 124.880 35.365 ;
        RECT 125.500 34.675 125.670 35.365 ;
        RECT 2.825 32.165 3.155 33.715 ;
        RECT 4.385 32.165 4.715 33.715 ;
        RECT 5.945 32.165 6.275 33.795 ;
        RECT 8.845 32.725 9.175 33.795 ;
        RECT 10.450 32.895 10.780 33.795 ;
        RECT 11.930 33.080 12.180 33.815 ;
        RECT 13.490 33.080 14.075 33.815 ;
        RECT 11.930 32.910 14.075 33.080 ;
        RECT 15.925 33.085 16.135 33.580 ;
        RECT 17.485 33.085 17.695 33.580 ;
        RECT 19.045 33.085 19.255 33.580 ;
        RECT 20.645 33.085 21.295 33.580 ;
        RECT 15.925 32.910 21.840 33.085 ;
        RECT 7.990 32.165 8.320 32.725 ;
        RECT 2.825 31.835 8.320 32.165 ;
        RECT 3.215 29.225 3.505 31.665 ;
        RECT 6.515 29.635 6.845 31.835 ;
        RECT 7.990 31.375 8.320 31.835 ;
        RECT 8.845 32.395 10.370 32.725 ;
        RECT 7.015 30.640 7.825 30.970 ;
        RECT 7.495 29.975 7.825 30.640 ;
        RECT 8.845 30.575 9.175 32.395 ;
        RECT 10.540 32.225 10.780 32.895 ;
        RECT 13.905 32.760 14.075 32.910 ;
        RECT 13.905 32.730 14.605 32.760 ;
        RECT 11.015 32.560 13.725 32.730 ;
        RECT 13.905 32.495 21.490 32.730 ;
        RECT 13.905 32.380 15.710 32.495 ;
        RECT 10.450 30.575 10.780 32.225 ;
        RECT 11.930 32.210 15.710 32.380 ;
        RECT 21.670 32.280 21.840 32.910 ;
        RECT 16.045 32.275 21.840 32.280 ;
        RECT 11.930 30.555 12.260 32.210 ;
        RECT 13.570 30.555 13.820 32.210 ;
        RECT 16.005 32.105 21.840 32.275 ;
        RECT 16.005 30.865 16.335 32.105 ;
        RECT 17.565 30.865 17.895 32.105 ;
        RECT 19.125 30.865 19.455 32.105 ;
        RECT 20.685 30.865 21.015 32.105 ;
        RECT 6.515 29.305 7.325 29.635 ;
        RECT 3.215 28.935 3.595 29.225 ;
        RECT 3.305 28.165 3.595 28.935 ;
        RECT 4.205 28.645 4.515 29.075 ;
        RECT 6.995 28.965 7.325 29.305 ;
        RECT 7.495 29.565 8.165 29.975 ;
        RECT 7.495 28.645 7.825 29.565 ;
        RECT 4.205 28.335 6.120 28.645 ;
        RECT 4.810 28.315 6.120 28.335 ;
        RECT 6.290 28.315 9.740 28.645 ;
        RECT 3.305 27.915 4.640 28.165 ;
        RECT 3.305 26.905 3.595 27.915 ;
        RECT 4.810 27.745 5.140 28.315 ;
        RECT 4.205 27.415 5.140 27.745 ;
        RECT 4.205 26.905 4.515 27.415 ;
        RECT 6.290 26.765 6.620 28.315 ;
        RECT 7.850 26.765 8.180 28.315 ;
        RECT 9.410 26.685 9.740 28.315 ;
        RECT 11.015 27.720 11.960 28.050 ;
        RECT 12.130 27.950 12.380 29.925 ;
        RECT 31.475 29.885 32.185 34.460 ;
        RECT 32.725 32.880 32.895 33.920 ;
        RECT 33.515 32.880 33.685 33.920 ;
        RECT 34.105 32.880 34.275 33.920 ;
        RECT 34.895 32.880 35.065 33.920 ;
        RECT 32.725 30.325 32.895 31.365 ;
        RECT 33.515 30.325 33.685 31.365 ;
        RECT 34.105 30.325 34.275 31.365 ;
        RECT 34.895 30.325 35.065 31.365 ;
        RECT 35.610 29.885 36.320 34.460 ;
        RECT 36.800 29.870 37.510 34.445 ;
        RECT 38.050 32.880 38.220 33.920 ;
        RECT 38.840 32.880 39.010 33.920 ;
        RECT 39.430 32.880 39.600 33.920 ;
        RECT 40.220 32.880 40.390 33.920 ;
        RECT 38.280 32.495 38.780 32.665 ;
        RECT 39.660 32.495 40.160 32.665 ;
        RECT 38.280 31.580 38.780 31.750 ;
        RECT 39.660 31.580 40.160 31.750 ;
        RECT 38.050 30.325 38.220 31.365 ;
        RECT 38.840 30.325 39.010 31.365 ;
        RECT 39.430 30.325 39.600 31.365 ;
        RECT 40.220 30.325 40.390 31.365 ;
        RECT 40.935 29.865 41.645 34.440 ;
        RECT 42.135 29.870 42.845 34.445 ;
        RECT 43.385 32.880 43.555 33.920 ;
        RECT 44.175 32.880 44.345 33.920 ;
        RECT 44.765 32.880 44.935 33.920 ;
        RECT 45.555 32.880 45.725 33.920 ;
        RECT 43.615 32.495 44.115 32.665 ;
        RECT 44.995 32.495 45.495 32.665 ;
        RECT 43.615 31.580 44.115 31.750 ;
        RECT 44.995 31.580 45.495 31.750 ;
        RECT 43.385 30.325 43.555 31.365 ;
        RECT 44.175 30.325 44.345 31.365 ;
        RECT 44.765 30.325 44.935 31.365 ;
        RECT 45.555 30.325 45.725 31.365 ;
        RECT 46.270 29.865 46.980 34.440 ;
        RECT 47.460 29.870 48.170 34.445 ;
        RECT 48.710 32.880 48.880 33.920 ;
        RECT 49.500 32.880 49.670 33.920 ;
        RECT 50.090 32.880 50.260 33.920 ;
        RECT 50.880 32.880 51.050 33.920 ;
        RECT 48.940 32.495 49.440 32.665 ;
        RECT 50.320 32.495 50.820 32.665 ;
        RECT 48.940 31.580 49.440 31.750 ;
        RECT 50.320 31.580 50.820 31.750 ;
        RECT 48.710 30.325 48.880 31.365 ;
        RECT 49.500 30.325 49.670 31.365 ;
        RECT 50.090 30.325 50.260 31.365 ;
        RECT 50.880 30.325 51.050 31.365 ;
        RECT 51.595 29.865 52.305 34.440 ;
        RECT 52.795 29.870 53.505 34.445 ;
        RECT 54.045 32.880 54.215 33.920 ;
        RECT 54.835 32.880 55.005 33.920 ;
        RECT 55.425 32.880 55.595 33.920 ;
        RECT 56.215 32.880 56.385 33.920 ;
        RECT 54.275 32.495 54.775 32.665 ;
        RECT 55.655 32.495 56.155 32.665 ;
        RECT 54.275 31.580 54.775 31.750 ;
        RECT 55.655 31.580 56.155 31.750 ;
        RECT 54.045 30.325 54.215 31.365 ;
        RECT 54.835 30.325 55.005 31.365 ;
        RECT 55.425 30.325 55.595 31.365 ;
        RECT 56.215 30.325 56.385 31.365 ;
        RECT 56.930 29.865 57.640 34.440 ;
        RECT 58.120 29.870 58.830 34.445 ;
        RECT 59.370 32.880 59.540 33.920 ;
        RECT 60.160 32.880 60.330 33.920 ;
        RECT 60.750 32.880 60.920 33.920 ;
        RECT 61.540 32.880 61.710 33.920 ;
        RECT 59.600 32.495 60.100 32.665 ;
        RECT 60.980 32.495 61.480 32.665 ;
        RECT 59.600 31.580 60.100 31.750 ;
        RECT 60.980 31.580 61.480 31.750 ;
        RECT 59.370 30.325 59.540 31.365 ;
        RECT 60.160 30.325 60.330 31.365 ;
        RECT 60.750 30.325 60.920 31.365 ;
        RECT 61.540 30.325 61.710 31.365 ;
        RECT 62.255 29.865 62.965 34.440 ;
        RECT 63.455 29.870 64.165 34.445 ;
        RECT 64.705 32.880 64.875 33.920 ;
        RECT 65.495 32.880 65.665 33.920 ;
        RECT 66.085 32.880 66.255 33.920 ;
        RECT 66.875 32.880 67.045 33.920 ;
        RECT 64.935 32.495 65.435 32.665 ;
        RECT 66.315 32.495 66.815 32.665 ;
        RECT 64.935 31.580 65.435 31.750 ;
        RECT 66.315 31.580 66.815 31.750 ;
        RECT 64.705 30.325 64.875 31.365 ;
        RECT 65.495 30.325 65.665 31.365 ;
        RECT 66.085 30.325 66.255 31.365 ;
        RECT 66.875 30.325 67.045 31.365 ;
        RECT 67.590 29.865 68.300 34.440 ;
        RECT 68.780 29.870 69.490 34.445 ;
        RECT 70.030 32.880 70.200 33.920 ;
        RECT 70.820 32.880 70.990 33.920 ;
        RECT 71.410 32.880 71.580 33.920 ;
        RECT 72.200 32.880 72.370 33.920 ;
        RECT 70.260 32.495 70.760 32.665 ;
        RECT 71.640 32.495 72.140 32.665 ;
        RECT 70.260 31.580 70.760 31.750 ;
        RECT 71.640 31.580 72.140 31.750 ;
        RECT 70.030 30.325 70.200 31.365 ;
        RECT 70.820 30.325 70.990 31.365 ;
        RECT 71.410 30.325 71.580 31.365 ;
        RECT 72.200 30.325 72.370 31.365 ;
        RECT 72.915 29.865 73.625 34.440 ;
        RECT 74.115 29.870 74.825 34.445 ;
        RECT 75.365 32.880 75.535 33.920 ;
        RECT 76.155 32.880 76.325 33.920 ;
        RECT 76.745 32.880 76.915 33.920 ;
        RECT 77.535 32.880 77.705 33.920 ;
        RECT 75.595 32.495 76.095 32.665 ;
        RECT 76.975 32.495 77.475 32.665 ;
        RECT 75.595 31.580 76.095 31.750 ;
        RECT 76.975 31.580 77.475 31.750 ;
        RECT 75.365 30.325 75.535 31.365 ;
        RECT 76.155 30.325 76.325 31.365 ;
        RECT 76.745 30.325 76.915 31.365 ;
        RECT 77.535 30.325 77.705 31.365 ;
        RECT 78.250 29.865 78.960 34.440 ;
        RECT 79.440 29.870 80.150 34.445 ;
        RECT 80.690 32.880 80.860 33.920 ;
        RECT 81.480 32.880 81.650 33.920 ;
        RECT 82.070 32.880 82.240 33.920 ;
        RECT 82.860 32.880 83.030 33.920 ;
        RECT 80.920 32.495 81.420 32.665 ;
        RECT 82.300 32.495 82.800 32.665 ;
        RECT 80.920 31.580 81.420 31.750 ;
        RECT 82.300 31.580 82.800 31.750 ;
        RECT 80.690 30.325 80.860 31.365 ;
        RECT 81.480 30.325 81.650 31.365 ;
        RECT 82.070 30.325 82.240 31.365 ;
        RECT 82.860 30.325 83.030 31.365 ;
        RECT 83.575 29.865 84.285 34.440 ;
        RECT 84.775 29.870 85.485 34.445 ;
        RECT 86.025 32.880 86.195 33.920 ;
        RECT 86.815 32.880 86.985 33.920 ;
        RECT 87.405 32.880 87.575 33.920 ;
        RECT 88.195 32.880 88.365 33.920 ;
        RECT 86.255 32.495 86.755 32.665 ;
        RECT 87.635 32.495 88.135 32.665 ;
        RECT 86.255 31.580 86.755 31.750 ;
        RECT 87.635 31.580 88.135 31.750 ;
        RECT 86.025 30.325 86.195 31.365 ;
        RECT 86.815 30.325 86.985 31.365 ;
        RECT 87.405 30.325 87.575 31.365 ;
        RECT 88.195 30.325 88.365 31.365 ;
        RECT 88.910 29.865 89.620 34.440 ;
        RECT 90.100 29.870 90.810 34.445 ;
        RECT 91.350 32.880 91.520 33.920 ;
        RECT 92.140 32.880 92.310 33.920 ;
        RECT 92.730 32.880 92.900 33.920 ;
        RECT 93.520 32.880 93.690 33.920 ;
        RECT 91.580 32.495 92.080 32.665 ;
        RECT 92.960 32.495 93.460 32.665 ;
        RECT 91.580 31.580 92.080 31.750 ;
        RECT 92.960 31.580 93.460 31.750 ;
        RECT 91.350 30.325 91.520 31.365 ;
        RECT 92.140 30.325 92.310 31.365 ;
        RECT 92.730 30.325 92.900 31.365 ;
        RECT 93.520 30.325 93.690 31.365 ;
        RECT 94.235 29.865 94.945 34.440 ;
        RECT 95.435 29.870 96.145 34.445 ;
        RECT 96.685 32.880 96.855 33.920 ;
        RECT 97.475 32.880 97.645 33.920 ;
        RECT 98.065 32.880 98.235 33.920 ;
        RECT 98.855 32.880 99.025 33.920 ;
        RECT 96.915 32.495 97.415 32.665 ;
        RECT 98.295 32.495 98.795 32.665 ;
        RECT 96.915 31.580 97.415 31.750 ;
        RECT 98.295 31.580 98.795 31.750 ;
        RECT 96.685 30.325 96.855 31.365 ;
        RECT 97.475 30.325 97.645 31.365 ;
        RECT 98.065 30.325 98.235 31.365 ;
        RECT 98.855 30.325 99.025 31.365 ;
        RECT 99.570 29.865 100.280 34.440 ;
        RECT 100.760 29.870 101.470 34.445 ;
        RECT 102.010 32.880 102.180 33.920 ;
        RECT 102.800 32.880 102.970 33.920 ;
        RECT 103.390 32.880 103.560 33.920 ;
        RECT 104.180 32.880 104.350 33.920 ;
        RECT 102.240 32.495 102.740 32.665 ;
        RECT 103.620 32.495 104.120 32.665 ;
        RECT 102.240 31.580 102.740 31.750 ;
        RECT 103.620 31.580 104.120 31.750 ;
        RECT 102.010 30.325 102.180 31.365 ;
        RECT 102.800 30.325 102.970 31.365 ;
        RECT 103.390 30.325 103.560 31.365 ;
        RECT 104.180 30.325 104.350 31.365 ;
        RECT 104.895 29.865 105.605 34.440 ;
        RECT 106.095 29.870 106.805 34.445 ;
        RECT 107.345 32.880 107.515 33.920 ;
        RECT 108.135 32.880 108.305 33.920 ;
        RECT 108.725 32.880 108.895 33.920 ;
        RECT 109.515 32.880 109.685 33.920 ;
        RECT 107.575 32.495 108.075 32.665 ;
        RECT 108.955 32.495 109.455 32.665 ;
        RECT 107.575 31.580 108.075 31.750 ;
        RECT 108.955 31.580 109.455 31.750 ;
        RECT 107.345 30.325 107.515 31.365 ;
        RECT 108.135 30.325 108.305 31.365 ;
        RECT 108.725 30.325 108.895 31.365 ;
        RECT 109.515 30.325 109.685 31.365 ;
        RECT 110.230 29.865 110.940 34.440 ;
        RECT 111.420 29.870 112.130 34.445 ;
        RECT 112.670 32.880 112.840 33.920 ;
        RECT 113.460 32.880 113.630 33.920 ;
        RECT 114.050 32.880 114.220 33.920 ;
        RECT 114.840 32.880 115.010 33.920 ;
        RECT 112.900 32.495 113.400 32.665 ;
        RECT 114.280 32.495 114.780 32.665 ;
        RECT 112.900 31.580 113.400 31.750 ;
        RECT 114.280 31.580 114.780 31.750 ;
        RECT 112.670 30.325 112.840 31.365 ;
        RECT 113.460 30.325 113.630 31.365 ;
        RECT 114.050 30.325 114.220 31.365 ;
        RECT 114.840 30.325 115.010 31.365 ;
        RECT 115.555 29.865 116.265 34.440 ;
        RECT 116.755 29.870 117.465 34.445 ;
        RECT 118.005 32.880 118.175 33.920 ;
        RECT 118.795 32.880 118.965 33.920 ;
        RECT 119.385 32.880 119.555 33.920 ;
        RECT 120.175 32.880 120.345 33.920 ;
        RECT 118.235 32.495 118.735 32.665 ;
        RECT 119.615 32.495 120.115 32.665 ;
        RECT 118.235 31.580 118.735 31.750 ;
        RECT 119.615 31.580 120.115 31.750 ;
        RECT 118.005 30.325 118.175 31.365 ;
        RECT 118.795 30.325 118.965 31.365 ;
        RECT 119.385 30.325 119.555 31.365 ;
        RECT 120.175 30.325 120.345 31.365 ;
        RECT 120.890 29.865 121.600 34.440 ;
        RECT 122.080 29.885 122.790 34.460 ;
        RECT 123.330 32.880 123.500 33.920 ;
        RECT 124.120 32.880 124.290 33.920 ;
        RECT 124.710 32.880 124.880 33.920 ;
        RECT 125.500 32.880 125.670 33.920 ;
        RECT 123.330 30.325 123.500 31.365 ;
        RECT 124.120 30.325 124.290 31.365 ;
        RECT 124.710 30.325 124.880 31.365 ;
        RECT 125.500 30.325 125.670 31.365 ;
        RECT 126.215 29.885 126.925 34.460 ;
        RECT 14.565 28.375 14.895 29.615 ;
        RECT 16.125 28.375 16.455 29.615 ;
        RECT 17.685 28.375 18.015 29.615 ;
        RECT 19.245 28.375 19.575 29.615 ;
        RECT 32.725 28.880 32.895 29.570 ;
        RECT 33.515 28.880 33.685 29.570 ;
        RECT 34.105 28.880 34.275 29.570 ;
        RECT 34.895 28.880 35.065 29.570 ;
        RECT 38.050 28.880 38.220 29.570 ;
        RECT 38.840 28.880 39.010 29.570 ;
        RECT 39.430 28.880 39.600 29.570 ;
        RECT 40.220 28.880 40.390 29.570 ;
        RECT 43.385 28.880 43.555 29.570 ;
        RECT 44.175 28.880 44.345 29.570 ;
        RECT 44.765 28.880 44.935 29.570 ;
        RECT 45.555 28.880 45.725 29.570 ;
        RECT 48.710 28.880 48.880 29.570 ;
        RECT 49.500 28.880 49.670 29.570 ;
        RECT 50.090 28.880 50.260 29.570 ;
        RECT 50.880 28.880 51.050 29.570 ;
        RECT 54.045 28.880 54.215 29.570 ;
        RECT 54.835 28.880 55.005 29.570 ;
        RECT 55.425 28.880 55.595 29.570 ;
        RECT 56.215 28.880 56.385 29.570 ;
        RECT 59.370 28.880 59.540 29.570 ;
        RECT 60.160 28.880 60.330 29.570 ;
        RECT 60.750 28.880 60.920 29.570 ;
        RECT 61.540 28.880 61.710 29.570 ;
        RECT 64.705 28.880 64.875 29.570 ;
        RECT 65.495 28.880 65.665 29.570 ;
        RECT 66.085 28.880 66.255 29.570 ;
        RECT 66.875 28.880 67.045 29.570 ;
        RECT 70.030 28.880 70.200 29.570 ;
        RECT 70.820 28.880 70.990 29.570 ;
        RECT 71.410 28.880 71.580 29.570 ;
        RECT 72.200 28.880 72.370 29.570 ;
        RECT 75.365 28.880 75.535 29.570 ;
        RECT 76.155 28.880 76.325 29.570 ;
        RECT 76.745 28.880 76.915 29.570 ;
        RECT 77.535 28.880 77.705 29.570 ;
        RECT 80.690 28.880 80.860 29.570 ;
        RECT 81.480 28.880 81.650 29.570 ;
        RECT 82.070 28.880 82.240 29.570 ;
        RECT 82.860 28.880 83.030 29.570 ;
        RECT 86.025 28.880 86.195 29.570 ;
        RECT 86.815 28.880 86.985 29.570 ;
        RECT 87.405 28.880 87.575 29.570 ;
        RECT 88.195 28.880 88.365 29.570 ;
        RECT 91.350 28.880 91.520 29.570 ;
        RECT 92.140 28.880 92.310 29.570 ;
        RECT 92.730 28.880 92.900 29.570 ;
        RECT 93.520 28.880 93.690 29.570 ;
        RECT 96.685 28.880 96.855 29.570 ;
        RECT 97.475 28.880 97.645 29.570 ;
        RECT 98.065 28.880 98.235 29.570 ;
        RECT 98.855 28.880 99.025 29.570 ;
        RECT 102.010 28.880 102.180 29.570 ;
        RECT 102.800 28.880 102.970 29.570 ;
        RECT 103.390 28.880 103.560 29.570 ;
        RECT 104.180 28.880 104.350 29.570 ;
        RECT 107.345 28.880 107.515 29.570 ;
        RECT 108.135 28.880 108.305 29.570 ;
        RECT 108.725 28.880 108.895 29.570 ;
        RECT 109.515 28.880 109.685 29.570 ;
        RECT 112.670 28.880 112.840 29.570 ;
        RECT 113.460 28.880 113.630 29.570 ;
        RECT 114.050 28.880 114.220 29.570 ;
        RECT 114.840 28.880 115.010 29.570 ;
        RECT 118.005 28.880 118.175 29.570 ;
        RECT 118.795 28.880 118.965 29.570 ;
        RECT 119.385 28.880 119.555 29.570 ;
        RECT 120.175 28.880 120.345 29.570 ;
        RECT 123.330 28.880 123.500 29.570 ;
        RECT 124.120 28.880 124.290 29.570 ;
        RECT 124.710 28.880 124.880 29.570 ;
        RECT 125.500 28.880 125.670 29.570 ;
        RECT 38.280 28.540 38.780 28.710 ;
        RECT 39.660 28.540 40.160 28.710 ;
        RECT 43.615 28.540 44.115 28.710 ;
        RECT 44.995 28.540 45.495 28.710 ;
        RECT 48.940 28.540 49.440 28.710 ;
        RECT 50.320 28.540 50.820 28.710 ;
        RECT 54.275 28.540 54.775 28.710 ;
        RECT 55.655 28.540 56.155 28.710 ;
        RECT 59.600 28.540 60.100 28.710 ;
        RECT 60.980 28.540 61.480 28.710 ;
        RECT 64.935 28.540 65.435 28.710 ;
        RECT 66.315 28.540 66.815 28.710 ;
        RECT 70.260 28.540 70.760 28.710 ;
        RECT 71.640 28.540 72.140 28.710 ;
        RECT 75.595 28.540 76.095 28.710 ;
        RECT 76.975 28.540 77.475 28.710 ;
        RECT 80.920 28.540 81.420 28.710 ;
        RECT 82.300 28.540 82.800 28.710 ;
        RECT 86.255 28.540 86.755 28.710 ;
        RECT 87.635 28.540 88.135 28.710 ;
        RECT 91.580 28.540 92.080 28.710 ;
        RECT 92.960 28.540 93.460 28.710 ;
        RECT 96.915 28.540 97.415 28.710 ;
        RECT 98.295 28.540 98.795 28.710 ;
        RECT 102.240 28.540 102.740 28.710 ;
        RECT 103.620 28.540 104.120 28.710 ;
        RECT 107.575 28.540 108.075 28.710 ;
        RECT 108.955 28.540 109.455 28.710 ;
        RECT 112.900 28.540 113.400 28.710 ;
        RECT 114.280 28.540 114.780 28.710 ;
        RECT 118.235 28.540 118.735 28.710 ;
        RECT 119.615 28.540 120.115 28.710 ;
        RECT 14.565 28.205 20.400 28.375 ;
        RECT 16.175 28.190 20.400 28.205 ;
        RECT 14.645 27.985 15.945 28.015 ;
        RECT 12.130 27.780 12.685 27.950 ;
        RECT 12.455 27.540 12.685 27.780 ;
        RECT 13.600 27.750 20.050 27.985 ;
        RECT 12.090 26.710 12.685 27.540 ;
        RECT 14.485 27.565 19.515 27.570 ;
        RECT 20.230 27.565 20.400 28.190 ;
        RECT 38.280 28.000 38.780 28.170 ;
        RECT 39.660 28.000 40.160 28.170 ;
        RECT 43.615 28.000 44.115 28.170 ;
        RECT 44.995 28.000 45.495 28.170 ;
        RECT 48.940 28.000 49.440 28.170 ;
        RECT 50.320 28.000 50.820 28.170 ;
        RECT 54.275 28.000 54.775 28.170 ;
        RECT 55.655 28.000 56.155 28.170 ;
        RECT 59.600 28.000 60.100 28.170 ;
        RECT 60.980 28.000 61.480 28.170 ;
        RECT 64.935 28.000 65.435 28.170 ;
        RECT 66.315 28.000 66.815 28.170 ;
        RECT 70.260 28.000 70.760 28.170 ;
        RECT 71.640 28.000 72.140 28.170 ;
        RECT 75.595 28.000 76.095 28.170 ;
        RECT 76.975 28.000 77.475 28.170 ;
        RECT 80.920 28.000 81.420 28.170 ;
        RECT 82.300 28.000 82.800 28.170 ;
        RECT 86.255 28.000 86.755 28.170 ;
        RECT 87.635 28.000 88.135 28.170 ;
        RECT 91.580 28.000 92.080 28.170 ;
        RECT 92.960 28.000 93.460 28.170 ;
        RECT 96.915 28.000 97.415 28.170 ;
        RECT 98.295 28.000 98.795 28.170 ;
        RECT 102.240 28.000 102.740 28.170 ;
        RECT 103.620 28.000 104.120 28.170 ;
        RECT 107.575 28.000 108.075 28.170 ;
        RECT 108.955 28.000 109.455 28.170 ;
        RECT 112.900 28.000 113.400 28.170 ;
        RECT 114.280 28.000 114.780 28.170 ;
        RECT 118.235 28.000 118.735 28.170 ;
        RECT 119.615 28.000 120.115 28.170 ;
        RECT 14.485 27.400 20.400 27.565 ;
        RECT 14.485 26.900 14.695 27.400 ;
        RECT 16.045 27.395 20.400 27.400 ;
        RECT 16.045 27.385 20.260 27.395 ;
        RECT 16.045 26.900 16.255 27.385 ;
        RECT 17.605 26.900 17.815 27.385 ;
        RECT 19.205 26.900 19.855 27.385 ;
        RECT 32.725 27.140 32.895 27.830 ;
        RECT 33.515 27.140 33.685 27.830 ;
        RECT 34.105 27.140 34.275 27.830 ;
        RECT 34.895 27.140 35.065 27.830 ;
        RECT 38.050 27.140 38.220 27.830 ;
        RECT 38.840 27.140 39.010 27.830 ;
        RECT 39.430 27.140 39.600 27.830 ;
        RECT 40.220 27.140 40.390 27.830 ;
        RECT 43.385 27.140 43.555 27.830 ;
        RECT 44.175 27.140 44.345 27.830 ;
        RECT 44.765 27.140 44.935 27.830 ;
        RECT 45.555 27.140 45.725 27.830 ;
        RECT 48.710 27.140 48.880 27.830 ;
        RECT 49.500 27.140 49.670 27.830 ;
        RECT 50.090 27.140 50.260 27.830 ;
        RECT 50.880 27.140 51.050 27.830 ;
        RECT 54.045 27.140 54.215 27.830 ;
        RECT 54.835 27.140 55.005 27.830 ;
        RECT 55.425 27.140 55.595 27.830 ;
        RECT 56.215 27.140 56.385 27.830 ;
        RECT 59.370 27.140 59.540 27.830 ;
        RECT 60.160 27.140 60.330 27.830 ;
        RECT 60.750 27.140 60.920 27.830 ;
        RECT 61.540 27.140 61.710 27.830 ;
        RECT 64.705 27.140 64.875 27.830 ;
        RECT 65.495 27.140 65.665 27.830 ;
        RECT 66.085 27.140 66.255 27.830 ;
        RECT 66.875 27.140 67.045 27.830 ;
        RECT 70.030 27.140 70.200 27.830 ;
        RECT 70.820 27.140 70.990 27.830 ;
        RECT 71.410 27.140 71.580 27.830 ;
        RECT 72.200 27.140 72.370 27.830 ;
        RECT 75.365 27.140 75.535 27.830 ;
        RECT 76.155 27.140 76.325 27.830 ;
        RECT 76.745 27.140 76.915 27.830 ;
        RECT 77.535 27.140 77.705 27.830 ;
        RECT 80.690 27.140 80.860 27.830 ;
        RECT 81.480 27.140 81.650 27.830 ;
        RECT 82.070 27.140 82.240 27.830 ;
        RECT 82.860 27.140 83.030 27.830 ;
        RECT 86.025 27.140 86.195 27.830 ;
        RECT 86.815 27.140 86.985 27.830 ;
        RECT 87.405 27.140 87.575 27.830 ;
        RECT 88.195 27.140 88.365 27.830 ;
        RECT 91.350 27.140 91.520 27.830 ;
        RECT 92.140 27.140 92.310 27.830 ;
        RECT 92.730 27.140 92.900 27.830 ;
        RECT 93.520 27.140 93.690 27.830 ;
        RECT 96.685 27.140 96.855 27.830 ;
        RECT 97.475 27.140 97.645 27.830 ;
        RECT 98.065 27.140 98.235 27.830 ;
        RECT 98.855 27.140 99.025 27.830 ;
        RECT 102.010 27.140 102.180 27.830 ;
        RECT 102.800 27.140 102.970 27.830 ;
        RECT 103.390 27.140 103.560 27.830 ;
        RECT 104.180 27.140 104.350 27.830 ;
        RECT 107.345 27.140 107.515 27.830 ;
        RECT 108.135 27.140 108.305 27.830 ;
        RECT 108.725 27.140 108.895 27.830 ;
        RECT 109.515 27.140 109.685 27.830 ;
        RECT 112.670 27.140 112.840 27.830 ;
        RECT 113.460 27.140 113.630 27.830 ;
        RECT 114.050 27.140 114.220 27.830 ;
        RECT 114.840 27.140 115.010 27.830 ;
        RECT 118.005 27.140 118.175 27.830 ;
        RECT 118.795 27.140 118.965 27.830 ;
        RECT 119.385 27.140 119.555 27.830 ;
        RECT 120.175 27.140 120.345 27.830 ;
        RECT 123.330 27.140 123.500 27.830 ;
        RECT 124.120 27.140 124.290 27.830 ;
        RECT 124.710 27.140 124.880 27.830 ;
        RECT 125.500 27.140 125.670 27.830 ;
        RECT 2.825 24.025 3.155 25.575 ;
        RECT 4.385 24.025 4.715 25.575 ;
        RECT 5.945 24.025 6.275 25.655 ;
        RECT 8.845 24.585 9.175 25.655 ;
        RECT 10.450 24.755 10.780 25.655 ;
        RECT 11.930 24.940 12.180 25.675 ;
        RECT 13.490 24.940 14.075 25.675 ;
        RECT 11.930 24.770 14.075 24.940 ;
        RECT 15.925 24.945 16.135 25.440 ;
        RECT 17.485 24.945 17.695 25.440 ;
        RECT 19.045 24.945 19.255 25.440 ;
        RECT 20.645 24.945 21.295 25.440 ;
        RECT 15.925 24.770 21.840 24.945 ;
        RECT 7.990 24.025 8.320 24.585 ;
        RECT 2.825 23.695 8.320 24.025 ;
        RECT 3.215 21.085 3.505 23.525 ;
        RECT 6.515 21.495 6.845 23.695 ;
        RECT 7.990 23.235 8.320 23.695 ;
        RECT 8.845 24.255 10.370 24.585 ;
        RECT 7.015 22.500 7.825 22.830 ;
        RECT 7.495 21.835 7.825 22.500 ;
        RECT 8.845 22.435 9.175 24.255 ;
        RECT 10.540 24.085 10.780 24.755 ;
        RECT 13.905 24.620 14.075 24.770 ;
        RECT 13.905 24.590 14.605 24.620 ;
        RECT 11.015 24.420 13.725 24.590 ;
        RECT 13.905 24.355 21.490 24.590 ;
        RECT 13.905 24.240 15.710 24.355 ;
        RECT 10.450 22.435 10.780 24.085 ;
        RECT 11.930 24.070 15.710 24.240 ;
        RECT 21.670 24.140 21.840 24.770 ;
        RECT 16.045 24.135 21.840 24.140 ;
        RECT 11.930 22.415 12.260 24.070 ;
        RECT 13.570 22.415 13.820 24.070 ;
        RECT 16.005 23.965 21.840 24.135 ;
        RECT 16.005 22.725 16.335 23.965 ;
        RECT 17.565 22.725 17.895 23.965 ;
        RECT 19.125 22.725 19.455 23.965 ;
        RECT 20.685 22.725 21.015 23.965 ;
        RECT 31.475 22.350 32.185 26.925 ;
        RECT 32.725 25.345 32.895 26.385 ;
        RECT 33.515 25.345 33.685 26.385 ;
        RECT 34.105 25.345 34.275 26.385 ;
        RECT 34.895 25.345 35.065 26.385 ;
        RECT 32.725 22.790 32.895 23.830 ;
        RECT 33.515 22.790 33.685 23.830 ;
        RECT 34.105 22.790 34.275 23.830 ;
        RECT 34.895 22.790 35.065 23.830 ;
        RECT 35.610 22.350 36.320 26.925 ;
        RECT 36.800 22.335 37.510 26.910 ;
        RECT 38.050 25.345 38.220 26.385 ;
        RECT 38.840 25.345 39.010 26.385 ;
        RECT 39.430 25.345 39.600 26.385 ;
        RECT 40.220 25.345 40.390 26.385 ;
        RECT 38.280 24.960 38.780 25.130 ;
        RECT 39.660 24.960 40.160 25.130 ;
        RECT 38.280 24.045 38.780 24.215 ;
        RECT 39.660 24.045 40.160 24.215 ;
        RECT 38.050 22.790 38.220 23.830 ;
        RECT 38.840 22.790 39.010 23.830 ;
        RECT 39.430 22.790 39.600 23.830 ;
        RECT 40.220 22.790 40.390 23.830 ;
        RECT 40.935 22.330 41.645 26.905 ;
        RECT 42.135 22.335 42.845 26.910 ;
        RECT 43.385 25.345 43.555 26.385 ;
        RECT 44.175 25.345 44.345 26.385 ;
        RECT 44.765 25.345 44.935 26.385 ;
        RECT 45.555 25.345 45.725 26.385 ;
        RECT 43.615 24.960 44.115 25.130 ;
        RECT 44.995 24.960 45.495 25.130 ;
        RECT 43.615 24.045 44.115 24.215 ;
        RECT 44.995 24.045 45.495 24.215 ;
        RECT 43.385 22.790 43.555 23.830 ;
        RECT 44.175 22.790 44.345 23.830 ;
        RECT 44.765 22.790 44.935 23.830 ;
        RECT 45.555 22.790 45.725 23.830 ;
        RECT 46.270 22.330 46.980 26.905 ;
        RECT 47.460 22.335 48.170 26.910 ;
        RECT 48.710 25.345 48.880 26.385 ;
        RECT 49.500 25.345 49.670 26.385 ;
        RECT 50.090 25.345 50.260 26.385 ;
        RECT 50.880 25.345 51.050 26.385 ;
        RECT 48.940 24.960 49.440 25.130 ;
        RECT 50.320 24.960 50.820 25.130 ;
        RECT 48.940 24.045 49.440 24.215 ;
        RECT 50.320 24.045 50.820 24.215 ;
        RECT 48.710 22.790 48.880 23.830 ;
        RECT 49.500 22.790 49.670 23.830 ;
        RECT 50.090 22.790 50.260 23.830 ;
        RECT 50.880 22.790 51.050 23.830 ;
        RECT 51.595 22.330 52.305 26.905 ;
        RECT 52.795 22.335 53.505 26.910 ;
        RECT 54.045 25.345 54.215 26.385 ;
        RECT 54.835 25.345 55.005 26.385 ;
        RECT 55.425 25.345 55.595 26.385 ;
        RECT 56.215 25.345 56.385 26.385 ;
        RECT 54.275 24.960 54.775 25.130 ;
        RECT 55.655 24.960 56.155 25.130 ;
        RECT 54.275 24.045 54.775 24.215 ;
        RECT 55.655 24.045 56.155 24.215 ;
        RECT 54.045 22.790 54.215 23.830 ;
        RECT 54.835 22.790 55.005 23.830 ;
        RECT 55.425 22.790 55.595 23.830 ;
        RECT 56.215 22.790 56.385 23.830 ;
        RECT 56.930 22.330 57.640 26.905 ;
        RECT 58.120 22.335 58.830 26.910 ;
        RECT 59.370 25.345 59.540 26.385 ;
        RECT 60.160 25.345 60.330 26.385 ;
        RECT 60.750 25.345 60.920 26.385 ;
        RECT 61.540 25.345 61.710 26.385 ;
        RECT 59.600 24.960 60.100 25.130 ;
        RECT 60.980 24.960 61.480 25.130 ;
        RECT 59.600 24.045 60.100 24.215 ;
        RECT 60.980 24.045 61.480 24.215 ;
        RECT 59.370 22.790 59.540 23.830 ;
        RECT 60.160 22.790 60.330 23.830 ;
        RECT 60.750 22.790 60.920 23.830 ;
        RECT 61.540 22.790 61.710 23.830 ;
        RECT 62.255 22.330 62.965 26.905 ;
        RECT 63.455 22.335 64.165 26.910 ;
        RECT 64.705 25.345 64.875 26.385 ;
        RECT 65.495 25.345 65.665 26.385 ;
        RECT 66.085 25.345 66.255 26.385 ;
        RECT 66.875 25.345 67.045 26.385 ;
        RECT 64.935 24.960 65.435 25.130 ;
        RECT 66.315 24.960 66.815 25.130 ;
        RECT 64.935 24.045 65.435 24.215 ;
        RECT 66.315 24.045 66.815 24.215 ;
        RECT 64.705 22.790 64.875 23.830 ;
        RECT 65.495 22.790 65.665 23.830 ;
        RECT 66.085 22.790 66.255 23.830 ;
        RECT 66.875 22.790 67.045 23.830 ;
        RECT 67.590 22.330 68.300 26.905 ;
        RECT 68.780 22.335 69.490 26.910 ;
        RECT 70.030 25.345 70.200 26.385 ;
        RECT 70.820 25.345 70.990 26.385 ;
        RECT 71.410 25.345 71.580 26.385 ;
        RECT 72.200 25.345 72.370 26.385 ;
        RECT 70.260 24.960 70.760 25.130 ;
        RECT 71.640 24.960 72.140 25.130 ;
        RECT 70.260 24.045 70.760 24.215 ;
        RECT 71.640 24.045 72.140 24.215 ;
        RECT 70.030 22.790 70.200 23.830 ;
        RECT 70.820 22.790 70.990 23.830 ;
        RECT 71.410 22.790 71.580 23.830 ;
        RECT 72.200 22.790 72.370 23.830 ;
        RECT 72.915 22.330 73.625 26.905 ;
        RECT 74.115 22.335 74.825 26.910 ;
        RECT 75.365 25.345 75.535 26.385 ;
        RECT 76.155 25.345 76.325 26.385 ;
        RECT 76.745 25.345 76.915 26.385 ;
        RECT 77.535 25.345 77.705 26.385 ;
        RECT 75.595 24.960 76.095 25.130 ;
        RECT 76.975 24.960 77.475 25.130 ;
        RECT 75.595 24.045 76.095 24.215 ;
        RECT 76.975 24.045 77.475 24.215 ;
        RECT 75.365 22.790 75.535 23.830 ;
        RECT 76.155 22.790 76.325 23.830 ;
        RECT 76.745 22.790 76.915 23.830 ;
        RECT 77.535 22.790 77.705 23.830 ;
        RECT 78.250 22.330 78.960 26.905 ;
        RECT 79.440 22.335 80.150 26.910 ;
        RECT 80.690 25.345 80.860 26.385 ;
        RECT 81.480 25.345 81.650 26.385 ;
        RECT 82.070 25.345 82.240 26.385 ;
        RECT 82.860 25.345 83.030 26.385 ;
        RECT 80.920 24.960 81.420 25.130 ;
        RECT 82.300 24.960 82.800 25.130 ;
        RECT 80.920 24.045 81.420 24.215 ;
        RECT 82.300 24.045 82.800 24.215 ;
        RECT 80.690 22.790 80.860 23.830 ;
        RECT 81.480 22.790 81.650 23.830 ;
        RECT 82.070 22.790 82.240 23.830 ;
        RECT 82.860 22.790 83.030 23.830 ;
        RECT 83.575 22.330 84.285 26.905 ;
        RECT 84.775 22.335 85.485 26.910 ;
        RECT 86.025 25.345 86.195 26.385 ;
        RECT 86.815 25.345 86.985 26.385 ;
        RECT 87.405 25.345 87.575 26.385 ;
        RECT 88.195 25.345 88.365 26.385 ;
        RECT 86.255 24.960 86.755 25.130 ;
        RECT 87.635 24.960 88.135 25.130 ;
        RECT 86.255 24.045 86.755 24.215 ;
        RECT 87.635 24.045 88.135 24.215 ;
        RECT 86.025 22.790 86.195 23.830 ;
        RECT 86.815 22.790 86.985 23.830 ;
        RECT 87.405 22.790 87.575 23.830 ;
        RECT 88.195 22.790 88.365 23.830 ;
        RECT 88.910 22.330 89.620 26.905 ;
        RECT 90.100 22.335 90.810 26.910 ;
        RECT 91.350 25.345 91.520 26.385 ;
        RECT 92.140 25.345 92.310 26.385 ;
        RECT 92.730 25.345 92.900 26.385 ;
        RECT 93.520 25.345 93.690 26.385 ;
        RECT 91.580 24.960 92.080 25.130 ;
        RECT 92.960 24.960 93.460 25.130 ;
        RECT 91.580 24.045 92.080 24.215 ;
        RECT 92.960 24.045 93.460 24.215 ;
        RECT 91.350 22.790 91.520 23.830 ;
        RECT 92.140 22.790 92.310 23.830 ;
        RECT 92.730 22.790 92.900 23.830 ;
        RECT 93.520 22.790 93.690 23.830 ;
        RECT 94.235 22.330 94.945 26.905 ;
        RECT 95.435 22.335 96.145 26.910 ;
        RECT 96.685 25.345 96.855 26.385 ;
        RECT 97.475 25.345 97.645 26.385 ;
        RECT 98.065 25.345 98.235 26.385 ;
        RECT 98.855 25.345 99.025 26.385 ;
        RECT 96.915 24.960 97.415 25.130 ;
        RECT 98.295 24.960 98.795 25.130 ;
        RECT 96.915 24.045 97.415 24.215 ;
        RECT 98.295 24.045 98.795 24.215 ;
        RECT 96.685 22.790 96.855 23.830 ;
        RECT 97.475 22.790 97.645 23.830 ;
        RECT 98.065 22.790 98.235 23.830 ;
        RECT 98.855 22.790 99.025 23.830 ;
        RECT 99.570 22.330 100.280 26.905 ;
        RECT 100.760 22.335 101.470 26.910 ;
        RECT 102.010 25.345 102.180 26.385 ;
        RECT 102.800 25.345 102.970 26.385 ;
        RECT 103.390 25.345 103.560 26.385 ;
        RECT 104.180 25.345 104.350 26.385 ;
        RECT 102.240 24.960 102.740 25.130 ;
        RECT 103.620 24.960 104.120 25.130 ;
        RECT 102.240 24.045 102.740 24.215 ;
        RECT 103.620 24.045 104.120 24.215 ;
        RECT 102.010 22.790 102.180 23.830 ;
        RECT 102.800 22.790 102.970 23.830 ;
        RECT 103.390 22.790 103.560 23.830 ;
        RECT 104.180 22.790 104.350 23.830 ;
        RECT 104.895 22.330 105.605 26.905 ;
        RECT 106.095 22.335 106.805 26.910 ;
        RECT 107.345 25.345 107.515 26.385 ;
        RECT 108.135 25.345 108.305 26.385 ;
        RECT 108.725 25.345 108.895 26.385 ;
        RECT 109.515 25.345 109.685 26.385 ;
        RECT 107.575 24.960 108.075 25.130 ;
        RECT 108.955 24.960 109.455 25.130 ;
        RECT 107.575 24.045 108.075 24.215 ;
        RECT 108.955 24.045 109.455 24.215 ;
        RECT 107.345 22.790 107.515 23.830 ;
        RECT 108.135 22.790 108.305 23.830 ;
        RECT 108.725 22.790 108.895 23.830 ;
        RECT 109.515 22.790 109.685 23.830 ;
        RECT 110.230 22.330 110.940 26.905 ;
        RECT 111.420 22.335 112.130 26.910 ;
        RECT 112.670 25.345 112.840 26.385 ;
        RECT 113.460 25.345 113.630 26.385 ;
        RECT 114.050 25.345 114.220 26.385 ;
        RECT 114.840 25.345 115.010 26.385 ;
        RECT 112.900 24.960 113.400 25.130 ;
        RECT 114.280 24.960 114.780 25.130 ;
        RECT 112.900 24.045 113.400 24.215 ;
        RECT 114.280 24.045 114.780 24.215 ;
        RECT 112.670 22.790 112.840 23.830 ;
        RECT 113.460 22.790 113.630 23.830 ;
        RECT 114.050 22.790 114.220 23.830 ;
        RECT 114.840 22.790 115.010 23.830 ;
        RECT 115.555 22.330 116.265 26.905 ;
        RECT 116.755 22.335 117.465 26.910 ;
        RECT 118.005 25.345 118.175 26.385 ;
        RECT 118.795 25.345 118.965 26.385 ;
        RECT 119.385 25.345 119.555 26.385 ;
        RECT 120.175 25.345 120.345 26.385 ;
        RECT 118.235 24.960 118.735 25.130 ;
        RECT 119.615 24.960 120.115 25.130 ;
        RECT 118.235 24.045 118.735 24.215 ;
        RECT 119.615 24.045 120.115 24.215 ;
        RECT 118.005 22.790 118.175 23.830 ;
        RECT 118.795 22.790 118.965 23.830 ;
        RECT 119.385 22.790 119.555 23.830 ;
        RECT 120.175 22.790 120.345 23.830 ;
        RECT 120.890 22.330 121.600 26.905 ;
        RECT 122.080 22.350 122.790 26.925 ;
        RECT 123.330 25.345 123.500 26.385 ;
        RECT 124.120 25.345 124.290 26.385 ;
        RECT 124.710 25.345 124.880 26.385 ;
        RECT 125.500 25.345 125.670 26.385 ;
        RECT 123.330 22.790 123.500 23.830 ;
        RECT 124.120 22.790 124.290 23.830 ;
        RECT 124.710 22.790 124.880 23.830 ;
        RECT 125.500 22.790 125.670 23.830 ;
        RECT 126.215 22.350 126.925 26.925 ;
        RECT 6.515 21.165 7.325 21.495 ;
        RECT 3.215 20.795 3.595 21.085 ;
        RECT 3.305 20.025 3.595 20.795 ;
        RECT 4.205 20.505 4.515 20.935 ;
        RECT 6.995 20.825 7.325 21.165 ;
        RECT 7.495 21.425 8.165 21.835 ;
        RECT 7.495 20.505 7.825 21.425 ;
        RECT 4.205 20.195 6.120 20.505 ;
        RECT 4.810 20.175 6.120 20.195 ;
        RECT 6.290 20.175 9.740 20.505 ;
        RECT 3.305 19.775 4.640 20.025 ;
        RECT 3.305 18.765 3.595 19.775 ;
        RECT 4.810 19.605 5.140 20.175 ;
        RECT 4.205 19.275 5.140 19.605 ;
        RECT 4.205 18.765 4.515 19.275 ;
        RECT 6.290 18.625 6.620 20.175 ;
        RECT 7.850 18.625 8.180 20.175 ;
        RECT 9.410 18.545 9.740 20.175 ;
        RECT 11.015 19.580 11.960 19.910 ;
        RECT 12.130 19.810 12.380 21.785 ;
        RECT 14.565 20.235 14.895 21.475 ;
        RECT 16.125 20.235 16.455 21.475 ;
        RECT 17.685 20.235 18.015 21.475 ;
        RECT 19.245 20.235 19.575 21.475 ;
        RECT 32.725 21.345 32.895 22.035 ;
        RECT 33.515 21.345 33.685 22.035 ;
        RECT 34.105 21.345 34.275 22.035 ;
        RECT 34.895 21.345 35.065 22.035 ;
        RECT 38.050 21.345 38.220 22.035 ;
        RECT 38.840 21.345 39.010 22.035 ;
        RECT 39.430 21.345 39.600 22.035 ;
        RECT 40.220 21.345 40.390 22.035 ;
        RECT 43.385 21.345 43.555 22.035 ;
        RECT 44.175 21.345 44.345 22.035 ;
        RECT 44.765 21.345 44.935 22.035 ;
        RECT 45.555 21.345 45.725 22.035 ;
        RECT 48.710 21.345 48.880 22.035 ;
        RECT 49.500 21.345 49.670 22.035 ;
        RECT 50.090 21.345 50.260 22.035 ;
        RECT 50.880 21.345 51.050 22.035 ;
        RECT 54.045 21.345 54.215 22.035 ;
        RECT 54.835 21.345 55.005 22.035 ;
        RECT 55.425 21.345 55.595 22.035 ;
        RECT 56.215 21.345 56.385 22.035 ;
        RECT 59.370 21.345 59.540 22.035 ;
        RECT 60.160 21.345 60.330 22.035 ;
        RECT 60.750 21.345 60.920 22.035 ;
        RECT 61.540 21.345 61.710 22.035 ;
        RECT 64.705 21.345 64.875 22.035 ;
        RECT 65.495 21.345 65.665 22.035 ;
        RECT 66.085 21.345 66.255 22.035 ;
        RECT 66.875 21.345 67.045 22.035 ;
        RECT 70.030 21.345 70.200 22.035 ;
        RECT 70.820 21.345 70.990 22.035 ;
        RECT 71.410 21.345 71.580 22.035 ;
        RECT 72.200 21.345 72.370 22.035 ;
        RECT 75.365 21.345 75.535 22.035 ;
        RECT 76.155 21.345 76.325 22.035 ;
        RECT 76.745 21.345 76.915 22.035 ;
        RECT 77.535 21.345 77.705 22.035 ;
        RECT 80.690 21.345 80.860 22.035 ;
        RECT 81.480 21.345 81.650 22.035 ;
        RECT 82.070 21.345 82.240 22.035 ;
        RECT 82.860 21.345 83.030 22.035 ;
        RECT 86.025 21.345 86.195 22.035 ;
        RECT 86.815 21.345 86.985 22.035 ;
        RECT 87.405 21.345 87.575 22.035 ;
        RECT 88.195 21.345 88.365 22.035 ;
        RECT 91.350 21.345 91.520 22.035 ;
        RECT 92.140 21.345 92.310 22.035 ;
        RECT 92.730 21.345 92.900 22.035 ;
        RECT 93.520 21.345 93.690 22.035 ;
        RECT 96.685 21.345 96.855 22.035 ;
        RECT 97.475 21.345 97.645 22.035 ;
        RECT 98.065 21.345 98.235 22.035 ;
        RECT 98.855 21.345 99.025 22.035 ;
        RECT 102.010 21.345 102.180 22.035 ;
        RECT 102.800 21.345 102.970 22.035 ;
        RECT 103.390 21.345 103.560 22.035 ;
        RECT 104.180 21.345 104.350 22.035 ;
        RECT 107.345 21.345 107.515 22.035 ;
        RECT 108.135 21.345 108.305 22.035 ;
        RECT 108.725 21.345 108.895 22.035 ;
        RECT 109.515 21.345 109.685 22.035 ;
        RECT 112.670 21.345 112.840 22.035 ;
        RECT 113.460 21.345 113.630 22.035 ;
        RECT 114.050 21.345 114.220 22.035 ;
        RECT 114.840 21.345 115.010 22.035 ;
        RECT 118.005 21.345 118.175 22.035 ;
        RECT 118.795 21.345 118.965 22.035 ;
        RECT 119.385 21.345 119.555 22.035 ;
        RECT 120.175 21.345 120.345 22.035 ;
        RECT 123.330 21.345 123.500 22.035 ;
        RECT 124.120 21.345 124.290 22.035 ;
        RECT 124.710 21.345 124.880 22.035 ;
        RECT 125.500 21.345 125.670 22.035 ;
        RECT 38.280 21.005 38.780 21.175 ;
        RECT 39.660 21.005 40.160 21.175 ;
        RECT 43.615 21.005 44.115 21.175 ;
        RECT 44.995 21.005 45.495 21.175 ;
        RECT 48.940 21.005 49.440 21.175 ;
        RECT 50.320 21.005 50.820 21.175 ;
        RECT 54.275 21.005 54.775 21.175 ;
        RECT 55.655 21.005 56.155 21.175 ;
        RECT 59.600 21.005 60.100 21.175 ;
        RECT 60.980 21.005 61.480 21.175 ;
        RECT 64.935 21.005 65.435 21.175 ;
        RECT 66.315 21.005 66.815 21.175 ;
        RECT 70.260 21.005 70.760 21.175 ;
        RECT 71.640 21.005 72.140 21.175 ;
        RECT 75.595 21.005 76.095 21.175 ;
        RECT 76.975 21.005 77.475 21.175 ;
        RECT 80.920 21.005 81.420 21.175 ;
        RECT 82.300 21.005 82.800 21.175 ;
        RECT 86.255 21.005 86.755 21.175 ;
        RECT 87.635 21.005 88.135 21.175 ;
        RECT 91.580 21.005 92.080 21.175 ;
        RECT 92.960 21.005 93.460 21.175 ;
        RECT 96.915 21.005 97.415 21.175 ;
        RECT 98.295 21.005 98.795 21.175 ;
        RECT 102.240 21.005 102.740 21.175 ;
        RECT 103.620 21.005 104.120 21.175 ;
        RECT 107.575 21.005 108.075 21.175 ;
        RECT 108.955 21.005 109.455 21.175 ;
        RECT 112.900 21.005 113.400 21.175 ;
        RECT 114.280 21.005 114.780 21.175 ;
        RECT 118.235 21.005 118.735 21.175 ;
        RECT 119.615 21.005 120.115 21.175 ;
        RECT 38.280 20.465 38.780 20.635 ;
        RECT 39.660 20.465 40.160 20.635 ;
        RECT 43.615 20.465 44.115 20.635 ;
        RECT 44.995 20.465 45.495 20.635 ;
        RECT 48.940 20.465 49.440 20.635 ;
        RECT 50.320 20.465 50.820 20.635 ;
        RECT 54.275 20.465 54.775 20.635 ;
        RECT 55.655 20.465 56.155 20.635 ;
        RECT 59.600 20.465 60.100 20.635 ;
        RECT 60.980 20.465 61.480 20.635 ;
        RECT 64.935 20.465 65.435 20.635 ;
        RECT 66.315 20.465 66.815 20.635 ;
        RECT 70.260 20.465 70.760 20.635 ;
        RECT 71.640 20.465 72.140 20.635 ;
        RECT 75.595 20.465 76.095 20.635 ;
        RECT 76.975 20.465 77.475 20.635 ;
        RECT 80.920 20.465 81.420 20.635 ;
        RECT 82.300 20.465 82.800 20.635 ;
        RECT 86.255 20.465 86.755 20.635 ;
        RECT 87.635 20.465 88.135 20.635 ;
        RECT 91.580 20.465 92.080 20.635 ;
        RECT 92.960 20.465 93.460 20.635 ;
        RECT 96.915 20.465 97.415 20.635 ;
        RECT 98.295 20.465 98.795 20.635 ;
        RECT 102.240 20.465 102.740 20.635 ;
        RECT 103.620 20.465 104.120 20.635 ;
        RECT 107.575 20.465 108.075 20.635 ;
        RECT 108.955 20.465 109.455 20.635 ;
        RECT 112.900 20.465 113.400 20.635 ;
        RECT 114.280 20.465 114.780 20.635 ;
        RECT 118.235 20.465 118.735 20.635 ;
        RECT 119.615 20.465 120.115 20.635 ;
        RECT 14.565 20.065 20.400 20.235 ;
        RECT 16.175 20.050 20.400 20.065 ;
        RECT 14.645 19.845 15.945 19.875 ;
        RECT 12.130 19.640 12.685 19.810 ;
        RECT 12.455 19.400 12.685 19.640 ;
        RECT 13.600 19.610 20.050 19.845 ;
        RECT 12.090 18.570 12.685 19.400 ;
        RECT 14.485 19.425 19.515 19.430 ;
        RECT 20.230 19.425 20.400 20.050 ;
        RECT 32.725 19.605 32.895 20.295 ;
        RECT 33.515 19.605 33.685 20.295 ;
        RECT 34.105 19.605 34.275 20.295 ;
        RECT 34.895 19.605 35.065 20.295 ;
        RECT 38.050 19.605 38.220 20.295 ;
        RECT 38.840 19.605 39.010 20.295 ;
        RECT 39.430 19.605 39.600 20.295 ;
        RECT 40.220 19.605 40.390 20.295 ;
        RECT 43.385 19.605 43.555 20.295 ;
        RECT 44.175 19.605 44.345 20.295 ;
        RECT 44.765 19.605 44.935 20.295 ;
        RECT 45.555 19.605 45.725 20.295 ;
        RECT 48.710 19.605 48.880 20.295 ;
        RECT 49.500 19.605 49.670 20.295 ;
        RECT 50.090 19.605 50.260 20.295 ;
        RECT 50.880 19.605 51.050 20.295 ;
        RECT 54.045 19.605 54.215 20.295 ;
        RECT 54.835 19.605 55.005 20.295 ;
        RECT 55.425 19.605 55.595 20.295 ;
        RECT 56.215 19.605 56.385 20.295 ;
        RECT 59.370 19.605 59.540 20.295 ;
        RECT 60.160 19.605 60.330 20.295 ;
        RECT 60.750 19.605 60.920 20.295 ;
        RECT 61.540 19.605 61.710 20.295 ;
        RECT 64.705 19.605 64.875 20.295 ;
        RECT 65.495 19.605 65.665 20.295 ;
        RECT 66.085 19.605 66.255 20.295 ;
        RECT 66.875 19.605 67.045 20.295 ;
        RECT 70.030 19.605 70.200 20.295 ;
        RECT 70.820 19.605 70.990 20.295 ;
        RECT 71.410 19.605 71.580 20.295 ;
        RECT 72.200 19.605 72.370 20.295 ;
        RECT 75.365 19.605 75.535 20.295 ;
        RECT 76.155 19.605 76.325 20.295 ;
        RECT 76.745 19.605 76.915 20.295 ;
        RECT 77.535 19.605 77.705 20.295 ;
        RECT 80.690 19.605 80.860 20.295 ;
        RECT 81.480 19.605 81.650 20.295 ;
        RECT 82.070 19.605 82.240 20.295 ;
        RECT 82.860 19.605 83.030 20.295 ;
        RECT 86.025 19.605 86.195 20.295 ;
        RECT 86.815 19.605 86.985 20.295 ;
        RECT 87.405 19.605 87.575 20.295 ;
        RECT 88.195 19.605 88.365 20.295 ;
        RECT 91.350 19.605 91.520 20.295 ;
        RECT 92.140 19.605 92.310 20.295 ;
        RECT 92.730 19.605 92.900 20.295 ;
        RECT 93.520 19.605 93.690 20.295 ;
        RECT 96.685 19.605 96.855 20.295 ;
        RECT 97.475 19.605 97.645 20.295 ;
        RECT 98.065 19.605 98.235 20.295 ;
        RECT 98.855 19.605 99.025 20.295 ;
        RECT 102.010 19.605 102.180 20.295 ;
        RECT 102.800 19.605 102.970 20.295 ;
        RECT 103.390 19.605 103.560 20.295 ;
        RECT 104.180 19.605 104.350 20.295 ;
        RECT 107.345 19.605 107.515 20.295 ;
        RECT 108.135 19.605 108.305 20.295 ;
        RECT 108.725 19.605 108.895 20.295 ;
        RECT 109.515 19.605 109.685 20.295 ;
        RECT 112.670 19.605 112.840 20.295 ;
        RECT 113.460 19.605 113.630 20.295 ;
        RECT 114.050 19.605 114.220 20.295 ;
        RECT 114.840 19.605 115.010 20.295 ;
        RECT 118.005 19.605 118.175 20.295 ;
        RECT 118.795 19.605 118.965 20.295 ;
        RECT 119.385 19.605 119.555 20.295 ;
        RECT 120.175 19.605 120.345 20.295 ;
        RECT 123.330 19.605 123.500 20.295 ;
        RECT 124.120 19.605 124.290 20.295 ;
        RECT 124.710 19.605 124.880 20.295 ;
        RECT 125.500 19.605 125.670 20.295 ;
        RECT 14.485 19.260 20.400 19.425 ;
        RECT 14.485 18.760 14.695 19.260 ;
        RECT 16.045 19.255 20.400 19.260 ;
        RECT 16.045 19.245 20.260 19.255 ;
        RECT 16.045 18.760 16.255 19.245 ;
        RECT 17.605 18.760 17.815 19.245 ;
        RECT 19.205 18.760 19.855 19.245 ;
        RECT 2.825 15.885 3.155 17.435 ;
        RECT 4.385 15.885 4.715 17.435 ;
        RECT 5.945 15.885 6.275 17.515 ;
        RECT 8.845 16.445 9.175 17.515 ;
        RECT 10.450 16.615 10.780 17.515 ;
        RECT 11.930 16.800 12.180 17.535 ;
        RECT 13.490 16.800 14.075 17.535 ;
        RECT 11.930 16.630 14.075 16.800 ;
        RECT 15.925 16.805 16.135 17.300 ;
        RECT 17.485 16.805 17.695 17.300 ;
        RECT 19.045 16.805 19.255 17.300 ;
        RECT 20.645 16.805 21.295 17.300 ;
        RECT 15.925 16.630 21.840 16.805 ;
        RECT 7.990 15.885 8.320 16.445 ;
        RECT 2.825 15.555 8.320 15.885 ;
        RECT 3.215 12.945 3.505 15.385 ;
        RECT 6.515 13.355 6.845 15.555 ;
        RECT 7.990 15.095 8.320 15.555 ;
        RECT 8.845 16.115 10.370 16.445 ;
        RECT 7.015 14.360 7.825 14.690 ;
        RECT 7.495 13.695 7.825 14.360 ;
        RECT 8.845 14.295 9.175 16.115 ;
        RECT 10.540 15.945 10.780 16.615 ;
        RECT 13.905 16.480 14.075 16.630 ;
        RECT 13.905 16.450 14.605 16.480 ;
        RECT 11.015 16.280 13.725 16.450 ;
        RECT 13.905 16.215 21.490 16.450 ;
        RECT 13.905 16.100 15.710 16.215 ;
        RECT 10.450 14.295 10.780 15.945 ;
        RECT 11.930 15.930 15.710 16.100 ;
        RECT 21.670 16.000 21.840 16.630 ;
        RECT 16.045 15.995 21.840 16.000 ;
        RECT 11.930 14.275 12.260 15.930 ;
        RECT 13.570 14.275 13.820 15.930 ;
        RECT 16.005 15.825 21.840 15.995 ;
        RECT 16.005 14.585 16.335 15.825 ;
        RECT 17.565 14.585 17.895 15.825 ;
        RECT 19.125 14.585 19.455 15.825 ;
        RECT 20.685 14.585 21.015 15.825 ;
        RECT 31.475 14.815 32.185 19.390 ;
        RECT 32.725 17.810 32.895 18.850 ;
        RECT 33.515 17.810 33.685 18.850 ;
        RECT 34.105 17.810 34.275 18.850 ;
        RECT 34.895 17.810 35.065 18.850 ;
        RECT 32.725 15.255 32.895 16.295 ;
        RECT 33.515 15.255 33.685 16.295 ;
        RECT 34.105 15.255 34.275 16.295 ;
        RECT 34.895 15.255 35.065 16.295 ;
        RECT 35.610 14.815 36.320 19.390 ;
        RECT 36.800 14.800 37.510 19.375 ;
        RECT 38.050 17.810 38.220 18.850 ;
        RECT 38.840 17.810 39.010 18.850 ;
        RECT 39.430 17.810 39.600 18.850 ;
        RECT 40.220 17.810 40.390 18.850 ;
        RECT 38.280 17.425 38.780 17.595 ;
        RECT 39.660 17.425 40.160 17.595 ;
        RECT 38.280 16.510 38.780 16.680 ;
        RECT 39.660 16.510 40.160 16.680 ;
        RECT 38.050 15.255 38.220 16.295 ;
        RECT 38.840 15.255 39.010 16.295 ;
        RECT 39.430 15.255 39.600 16.295 ;
        RECT 40.220 15.255 40.390 16.295 ;
        RECT 40.935 14.795 41.645 19.370 ;
        RECT 42.135 14.800 42.845 19.375 ;
        RECT 43.385 17.810 43.555 18.850 ;
        RECT 44.175 17.810 44.345 18.850 ;
        RECT 44.765 17.810 44.935 18.850 ;
        RECT 45.555 17.810 45.725 18.850 ;
        RECT 43.615 17.425 44.115 17.595 ;
        RECT 44.995 17.425 45.495 17.595 ;
        RECT 43.615 16.510 44.115 16.680 ;
        RECT 44.995 16.510 45.495 16.680 ;
        RECT 43.385 15.255 43.555 16.295 ;
        RECT 44.175 15.255 44.345 16.295 ;
        RECT 44.765 15.255 44.935 16.295 ;
        RECT 45.555 15.255 45.725 16.295 ;
        RECT 46.270 14.795 46.980 19.370 ;
        RECT 47.460 14.800 48.170 19.375 ;
        RECT 48.710 17.810 48.880 18.850 ;
        RECT 49.500 17.810 49.670 18.850 ;
        RECT 50.090 17.810 50.260 18.850 ;
        RECT 50.880 17.810 51.050 18.850 ;
        RECT 48.940 17.425 49.440 17.595 ;
        RECT 50.320 17.425 50.820 17.595 ;
        RECT 48.940 16.510 49.440 16.680 ;
        RECT 50.320 16.510 50.820 16.680 ;
        RECT 48.710 15.255 48.880 16.295 ;
        RECT 49.500 15.255 49.670 16.295 ;
        RECT 50.090 15.255 50.260 16.295 ;
        RECT 50.880 15.255 51.050 16.295 ;
        RECT 51.595 14.795 52.305 19.370 ;
        RECT 52.795 14.800 53.505 19.375 ;
        RECT 54.045 17.810 54.215 18.850 ;
        RECT 54.835 17.810 55.005 18.850 ;
        RECT 55.425 17.810 55.595 18.850 ;
        RECT 56.215 17.810 56.385 18.850 ;
        RECT 54.275 17.425 54.775 17.595 ;
        RECT 55.655 17.425 56.155 17.595 ;
        RECT 54.275 16.510 54.775 16.680 ;
        RECT 55.655 16.510 56.155 16.680 ;
        RECT 54.045 15.255 54.215 16.295 ;
        RECT 54.835 15.255 55.005 16.295 ;
        RECT 55.425 15.255 55.595 16.295 ;
        RECT 56.215 15.255 56.385 16.295 ;
        RECT 56.930 14.795 57.640 19.370 ;
        RECT 58.120 14.800 58.830 19.375 ;
        RECT 59.370 17.810 59.540 18.850 ;
        RECT 60.160 17.810 60.330 18.850 ;
        RECT 60.750 17.810 60.920 18.850 ;
        RECT 61.540 17.810 61.710 18.850 ;
        RECT 59.600 17.425 60.100 17.595 ;
        RECT 60.980 17.425 61.480 17.595 ;
        RECT 59.600 16.510 60.100 16.680 ;
        RECT 60.980 16.510 61.480 16.680 ;
        RECT 59.370 15.255 59.540 16.295 ;
        RECT 60.160 15.255 60.330 16.295 ;
        RECT 60.750 15.255 60.920 16.295 ;
        RECT 61.540 15.255 61.710 16.295 ;
        RECT 62.255 14.795 62.965 19.370 ;
        RECT 63.455 14.800 64.165 19.375 ;
        RECT 64.705 17.810 64.875 18.850 ;
        RECT 65.495 17.810 65.665 18.850 ;
        RECT 66.085 17.810 66.255 18.850 ;
        RECT 66.875 17.810 67.045 18.850 ;
        RECT 64.935 17.425 65.435 17.595 ;
        RECT 66.315 17.425 66.815 17.595 ;
        RECT 64.935 16.510 65.435 16.680 ;
        RECT 66.315 16.510 66.815 16.680 ;
        RECT 64.705 15.255 64.875 16.295 ;
        RECT 65.495 15.255 65.665 16.295 ;
        RECT 66.085 15.255 66.255 16.295 ;
        RECT 66.875 15.255 67.045 16.295 ;
        RECT 67.590 14.795 68.300 19.370 ;
        RECT 68.780 14.800 69.490 19.375 ;
        RECT 70.030 17.810 70.200 18.850 ;
        RECT 70.820 17.810 70.990 18.850 ;
        RECT 71.410 17.810 71.580 18.850 ;
        RECT 72.200 17.810 72.370 18.850 ;
        RECT 70.260 17.425 70.760 17.595 ;
        RECT 71.640 17.425 72.140 17.595 ;
        RECT 70.260 16.510 70.760 16.680 ;
        RECT 71.640 16.510 72.140 16.680 ;
        RECT 70.030 15.255 70.200 16.295 ;
        RECT 70.820 15.255 70.990 16.295 ;
        RECT 71.410 15.255 71.580 16.295 ;
        RECT 72.200 15.255 72.370 16.295 ;
        RECT 72.915 14.795 73.625 19.370 ;
        RECT 74.115 14.800 74.825 19.375 ;
        RECT 75.365 17.810 75.535 18.850 ;
        RECT 76.155 17.810 76.325 18.850 ;
        RECT 76.745 17.810 76.915 18.850 ;
        RECT 77.535 17.810 77.705 18.850 ;
        RECT 75.595 17.425 76.095 17.595 ;
        RECT 76.975 17.425 77.475 17.595 ;
        RECT 75.595 16.510 76.095 16.680 ;
        RECT 76.975 16.510 77.475 16.680 ;
        RECT 75.365 15.255 75.535 16.295 ;
        RECT 76.155 15.255 76.325 16.295 ;
        RECT 76.745 15.255 76.915 16.295 ;
        RECT 77.535 15.255 77.705 16.295 ;
        RECT 78.250 14.795 78.960 19.370 ;
        RECT 79.440 14.800 80.150 19.375 ;
        RECT 80.690 17.810 80.860 18.850 ;
        RECT 81.480 17.810 81.650 18.850 ;
        RECT 82.070 17.810 82.240 18.850 ;
        RECT 82.860 17.810 83.030 18.850 ;
        RECT 80.920 17.425 81.420 17.595 ;
        RECT 82.300 17.425 82.800 17.595 ;
        RECT 80.920 16.510 81.420 16.680 ;
        RECT 82.300 16.510 82.800 16.680 ;
        RECT 80.690 15.255 80.860 16.295 ;
        RECT 81.480 15.255 81.650 16.295 ;
        RECT 82.070 15.255 82.240 16.295 ;
        RECT 82.860 15.255 83.030 16.295 ;
        RECT 83.575 14.795 84.285 19.370 ;
        RECT 84.775 14.800 85.485 19.375 ;
        RECT 86.025 17.810 86.195 18.850 ;
        RECT 86.815 17.810 86.985 18.850 ;
        RECT 87.405 17.810 87.575 18.850 ;
        RECT 88.195 17.810 88.365 18.850 ;
        RECT 86.255 17.425 86.755 17.595 ;
        RECT 87.635 17.425 88.135 17.595 ;
        RECT 86.255 16.510 86.755 16.680 ;
        RECT 87.635 16.510 88.135 16.680 ;
        RECT 86.025 15.255 86.195 16.295 ;
        RECT 86.815 15.255 86.985 16.295 ;
        RECT 87.405 15.255 87.575 16.295 ;
        RECT 88.195 15.255 88.365 16.295 ;
        RECT 88.910 14.795 89.620 19.370 ;
        RECT 90.100 14.800 90.810 19.375 ;
        RECT 91.350 17.810 91.520 18.850 ;
        RECT 92.140 17.810 92.310 18.850 ;
        RECT 92.730 17.810 92.900 18.850 ;
        RECT 93.520 17.810 93.690 18.850 ;
        RECT 91.580 17.425 92.080 17.595 ;
        RECT 92.960 17.425 93.460 17.595 ;
        RECT 91.580 16.510 92.080 16.680 ;
        RECT 92.960 16.510 93.460 16.680 ;
        RECT 91.350 15.255 91.520 16.295 ;
        RECT 92.140 15.255 92.310 16.295 ;
        RECT 92.730 15.255 92.900 16.295 ;
        RECT 93.520 15.255 93.690 16.295 ;
        RECT 94.235 14.795 94.945 19.370 ;
        RECT 95.435 14.800 96.145 19.375 ;
        RECT 96.685 17.810 96.855 18.850 ;
        RECT 97.475 17.810 97.645 18.850 ;
        RECT 98.065 17.810 98.235 18.850 ;
        RECT 98.855 17.810 99.025 18.850 ;
        RECT 96.915 17.425 97.415 17.595 ;
        RECT 98.295 17.425 98.795 17.595 ;
        RECT 96.915 16.510 97.415 16.680 ;
        RECT 98.295 16.510 98.795 16.680 ;
        RECT 96.685 15.255 96.855 16.295 ;
        RECT 97.475 15.255 97.645 16.295 ;
        RECT 98.065 15.255 98.235 16.295 ;
        RECT 98.855 15.255 99.025 16.295 ;
        RECT 99.570 14.795 100.280 19.370 ;
        RECT 100.760 14.800 101.470 19.375 ;
        RECT 102.010 17.810 102.180 18.850 ;
        RECT 102.800 17.810 102.970 18.850 ;
        RECT 103.390 17.810 103.560 18.850 ;
        RECT 104.180 17.810 104.350 18.850 ;
        RECT 102.240 17.425 102.740 17.595 ;
        RECT 103.620 17.425 104.120 17.595 ;
        RECT 102.240 16.510 102.740 16.680 ;
        RECT 103.620 16.510 104.120 16.680 ;
        RECT 102.010 15.255 102.180 16.295 ;
        RECT 102.800 15.255 102.970 16.295 ;
        RECT 103.390 15.255 103.560 16.295 ;
        RECT 104.180 15.255 104.350 16.295 ;
        RECT 104.895 14.795 105.605 19.370 ;
        RECT 106.095 14.800 106.805 19.375 ;
        RECT 107.345 17.810 107.515 18.850 ;
        RECT 108.135 17.810 108.305 18.850 ;
        RECT 108.725 17.810 108.895 18.850 ;
        RECT 109.515 17.810 109.685 18.850 ;
        RECT 107.575 17.425 108.075 17.595 ;
        RECT 108.955 17.425 109.455 17.595 ;
        RECT 107.575 16.510 108.075 16.680 ;
        RECT 108.955 16.510 109.455 16.680 ;
        RECT 107.345 15.255 107.515 16.295 ;
        RECT 108.135 15.255 108.305 16.295 ;
        RECT 108.725 15.255 108.895 16.295 ;
        RECT 109.515 15.255 109.685 16.295 ;
        RECT 110.230 14.795 110.940 19.370 ;
        RECT 111.420 14.800 112.130 19.375 ;
        RECT 112.670 17.810 112.840 18.850 ;
        RECT 113.460 17.810 113.630 18.850 ;
        RECT 114.050 17.810 114.220 18.850 ;
        RECT 114.840 17.810 115.010 18.850 ;
        RECT 112.900 17.425 113.400 17.595 ;
        RECT 114.280 17.425 114.780 17.595 ;
        RECT 112.900 16.510 113.400 16.680 ;
        RECT 114.280 16.510 114.780 16.680 ;
        RECT 112.670 15.255 112.840 16.295 ;
        RECT 113.460 15.255 113.630 16.295 ;
        RECT 114.050 15.255 114.220 16.295 ;
        RECT 114.840 15.255 115.010 16.295 ;
        RECT 115.555 14.795 116.265 19.370 ;
        RECT 116.755 14.800 117.465 19.375 ;
        RECT 118.005 17.810 118.175 18.850 ;
        RECT 118.795 17.810 118.965 18.850 ;
        RECT 119.385 17.810 119.555 18.850 ;
        RECT 120.175 17.810 120.345 18.850 ;
        RECT 118.235 17.425 118.735 17.595 ;
        RECT 119.615 17.425 120.115 17.595 ;
        RECT 118.235 16.510 118.735 16.680 ;
        RECT 119.615 16.510 120.115 16.680 ;
        RECT 118.005 15.255 118.175 16.295 ;
        RECT 118.795 15.255 118.965 16.295 ;
        RECT 119.385 15.255 119.555 16.295 ;
        RECT 120.175 15.255 120.345 16.295 ;
        RECT 120.890 14.795 121.600 19.370 ;
        RECT 122.080 14.815 122.790 19.390 ;
        RECT 123.330 17.810 123.500 18.850 ;
        RECT 124.120 17.810 124.290 18.850 ;
        RECT 124.710 17.810 124.880 18.850 ;
        RECT 125.500 17.810 125.670 18.850 ;
        RECT 123.330 15.255 123.500 16.295 ;
        RECT 124.120 15.255 124.290 16.295 ;
        RECT 124.710 15.255 124.880 16.295 ;
        RECT 125.500 15.255 125.670 16.295 ;
        RECT 126.215 14.815 126.925 19.390 ;
        RECT 32.725 13.810 32.895 14.500 ;
        RECT 33.515 13.810 33.685 14.500 ;
        RECT 34.105 13.810 34.275 14.500 ;
        RECT 34.895 13.810 35.065 14.500 ;
        RECT 38.050 13.810 38.220 14.500 ;
        RECT 38.840 13.810 39.010 14.500 ;
        RECT 39.430 13.810 39.600 14.500 ;
        RECT 40.220 13.810 40.390 14.500 ;
        RECT 43.385 13.810 43.555 14.500 ;
        RECT 44.175 13.810 44.345 14.500 ;
        RECT 44.765 13.810 44.935 14.500 ;
        RECT 45.555 13.810 45.725 14.500 ;
        RECT 48.710 13.810 48.880 14.500 ;
        RECT 49.500 13.810 49.670 14.500 ;
        RECT 50.090 13.810 50.260 14.500 ;
        RECT 50.880 13.810 51.050 14.500 ;
        RECT 54.045 13.810 54.215 14.500 ;
        RECT 54.835 13.810 55.005 14.500 ;
        RECT 55.425 13.810 55.595 14.500 ;
        RECT 56.215 13.810 56.385 14.500 ;
        RECT 59.370 13.810 59.540 14.500 ;
        RECT 60.160 13.810 60.330 14.500 ;
        RECT 60.750 13.810 60.920 14.500 ;
        RECT 61.540 13.810 61.710 14.500 ;
        RECT 64.705 13.810 64.875 14.500 ;
        RECT 65.495 13.810 65.665 14.500 ;
        RECT 66.085 13.810 66.255 14.500 ;
        RECT 66.875 13.810 67.045 14.500 ;
        RECT 70.030 13.810 70.200 14.500 ;
        RECT 70.820 13.810 70.990 14.500 ;
        RECT 71.410 13.810 71.580 14.500 ;
        RECT 72.200 13.810 72.370 14.500 ;
        RECT 75.365 13.810 75.535 14.500 ;
        RECT 76.155 13.810 76.325 14.500 ;
        RECT 76.745 13.810 76.915 14.500 ;
        RECT 77.535 13.810 77.705 14.500 ;
        RECT 80.690 13.810 80.860 14.500 ;
        RECT 81.480 13.810 81.650 14.500 ;
        RECT 82.070 13.810 82.240 14.500 ;
        RECT 82.860 13.810 83.030 14.500 ;
        RECT 86.025 13.810 86.195 14.500 ;
        RECT 86.815 13.810 86.985 14.500 ;
        RECT 87.405 13.810 87.575 14.500 ;
        RECT 88.195 13.810 88.365 14.500 ;
        RECT 91.350 13.810 91.520 14.500 ;
        RECT 92.140 13.810 92.310 14.500 ;
        RECT 92.730 13.810 92.900 14.500 ;
        RECT 93.520 13.810 93.690 14.500 ;
        RECT 96.685 13.810 96.855 14.500 ;
        RECT 97.475 13.810 97.645 14.500 ;
        RECT 98.065 13.810 98.235 14.500 ;
        RECT 98.855 13.810 99.025 14.500 ;
        RECT 102.010 13.810 102.180 14.500 ;
        RECT 102.800 13.810 102.970 14.500 ;
        RECT 103.390 13.810 103.560 14.500 ;
        RECT 104.180 13.810 104.350 14.500 ;
        RECT 107.345 13.810 107.515 14.500 ;
        RECT 108.135 13.810 108.305 14.500 ;
        RECT 108.725 13.810 108.895 14.500 ;
        RECT 109.515 13.810 109.685 14.500 ;
        RECT 112.670 13.810 112.840 14.500 ;
        RECT 113.460 13.810 113.630 14.500 ;
        RECT 114.050 13.810 114.220 14.500 ;
        RECT 114.840 13.810 115.010 14.500 ;
        RECT 118.005 13.810 118.175 14.500 ;
        RECT 118.795 13.810 118.965 14.500 ;
        RECT 119.385 13.810 119.555 14.500 ;
        RECT 120.175 13.810 120.345 14.500 ;
        RECT 123.330 13.810 123.500 14.500 ;
        RECT 124.120 13.810 124.290 14.500 ;
        RECT 124.710 13.810 124.880 14.500 ;
        RECT 125.500 13.810 125.670 14.500 ;
        RECT 6.515 13.025 7.325 13.355 ;
        RECT 3.215 12.655 3.595 12.945 ;
        RECT 3.305 11.885 3.595 12.655 ;
        RECT 4.205 12.365 4.515 12.795 ;
        RECT 6.995 12.685 7.325 13.025 ;
        RECT 7.495 13.285 8.165 13.695 ;
        RECT 7.495 12.365 7.825 13.285 ;
        RECT 4.205 12.055 6.120 12.365 ;
        RECT 4.810 12.035 6.120 12.055 ;
        RECT 6.290 12.035 9.740 12.365 ;
        RECT 3.305 11.635 4.640 11.885 ;
        RECT 3.305 10.625 3.595 11.635 ;
        RECT 4.810 11.465 5.140 12.035 ;
        RECT 4.205 11.135 5.140 11.465 ;
        RECT 4.205 10.625 4.515 11.135 ;
        RECT 6.290 10.485 6.620 12.035 ;
        RECT 7.850 10.485 8.180 12.035 ;
        RECT 9.410 10.405 9.740 12.035 ;
        RECT 11.015 11.440 11.960 11.770 ;
        RECT 12.130 11.670 12.380 13.645 ;
        RECT 38.280 13.470 38.780 13.640 ;
        RECT 39.660 13.470 40.160 13.640 ;
        RECT 43.615 13.470 44.115 13.640 ;
        RECT 44.995 13.470 45.495 13.640 ;
        RECT 48.940 13.470 49.440 13.640 ;
        RECT 50.320 13.470 50.820 13.640 ;
        RECT 54.275 13.470 54.775 13.640 ;
        RECT 55.655 13.470 56.155 13.640 ;
        RECT 59.600 13.470 60.100 13.640 ;
        RECT 60.980 13.470 61.480 13.640 ;
        RECT 64.935 13.470 65.435 13.640 ;
        RECT 66.315 13.470 66.815 13.640 ;
        RECT 70.260 13.470 70.760 13.640 ;
        RECT 71.640 13.470 72.140 13.640 ;
        RECT 75.595 13.470 76.095 13.640 ;
        RECT 76.975 13.470 77.475 13.640 ;
        RECT 80.920 13.470 81.420 13.640 ;
        RECT 82.300 13.470 82.800 13.640 ;
        RECT 86.255 13.470 86.755 13.640 ;
        RECT 87.635 13.470 88.135 13.640 ;
        RECT 91.580 13.470 92.080 13.640 ;
        RECT 92.960 13.470 93.460 13.640 ;
        RECT 96.915 13.470 97.415 13.640 ;
        RECT 98.295 13.470 98.795 13.640 ;
        RECT 102.240 13.470 102.740 13.640 ;
        RECT 103.620 13.470 104.120 13.640 ;
        RECT 107.575 13.470 108.075 13.640 ;
        RECT 108.955 13.470 109.455 13.640 ;
        RECT 112.900 13.470 113.400 13.640 ;
        RECT 114.280 13.470 114.780 13.640 ;
        RECT 118.235 13.470 118.735 13.640 ;
        RECT 119.615 13.470 120.115 13.640 ;
        RECT 14.565 12.095 14.895 13.335 ;
        RECT 16.125 12.095 16.455 13.335 ;
        RECT 17.685 12.095 18.015 13.335 ;
        RECT 19.245 12.095 19.575 13.335 ;
        RECT 38.280 12.930 38.780 13.100 ;
        RECT 39.660 12.930 40.160 13.100 ;
        RECT 43.615 12.930 44.115 13.100 ;
        RECT 44.995 12.930 45.495 13.100 ;
        RECT 48.940 12.930 49.440 13.100 ;
        RECT 50.320 12.930 50.820 13.100 ;
        RECT 54.275 12.930 54.775 13.100 ;
        RECT 55.655 12.930 56.155 13.100 ;
        RECT 59.600 12.930 60.100 13.100 ;
        RECT 60.980 12.930 61.480 13.100 ;
        RECT 64.935 12.930 65.435 13.100 ;
        RECT 66.315 12.930 66.815 13.100 ;
        RECT 70.260 12.930 70.760 13.100 ;
        RECT 71.640 12.930 72.140 13.100 ;
        RECT 75.595 12.930 76.095 13.100 ;
        RECT 76.975 12.930 77.475 13.100 ;
        RECT 80.920 12.930 81.420 13.100 ;
        RECT 82.300 12.930 82.800 13.100 ;
        RECT 86.255 12.930 86.755 13.100 ;
        RECT 87.635 12.930 88.135 13.100 ;
        RECT 91.580 12.930 92.080 13.100 ;
        RECT 92.960 12.930 93.460 13.100 ;
        RECT 96.915 12.930 97.415 13.100 ;
        RECT 98.295 12.930 98.795 13.100 ;
        RECT 102.240 12.930 102.740 13.100 ;
        RECT 103.620 12.930 104.120 13.100 ;
        RECT 107.575 12.930 108.075 13.100 ;
        RECT 108.955 12.930 109.455 13.100 ;
        RECT 112.900 12.930 113.400 13.100 ;
        RECT 114.280 12.930 114.780 13.100 ;
        RECT 118.235 12.930 118.735 13.100 ;
        RECT 119.615 12.930 120.115 13.100 ;
        RECT 14.565 11.925 20.400 12.095 ;
        RECT 32.725 12.070 32.895 12.760 ;
        RECT 33.515 12.070 33.685 12.760 ;
        RECT 34.105 12.070 34.275 12.760 ;
        RECT 34.895 12.070 35.065 12.760 ;
        RECT 38.840 12.070 39.010 12.760 ;
        RECT 39.430 12.070 39.600 12.760 ;
        RECT 40.220 12.070 40.390 12.760 ;
        RECT 43.385 12.070 43.555 12.760 ;
        RECT 44.175 12.070 44.345 12.760 ;
        RECT 44.765 12.070 44.935 12.760 ;
        RECT 45.555 12.070 45.725 12.760 ;
        RECT 48.710 12.070 48.880 12.760 ;
        RECT 49.500 12.070 49.670 12.760 ;
        RECT 50.090 12.070 50.260 12.760 ;
        RECT 50.880 12.070 51.050 12.760 ;
        RECT 54.045 12.070 54.215 12.760 ;
        RECT 54.835 12.070 55.005 12.760 ;
        RECT 55.425 12.070 55.595 12.760 ;
        RECT 56.215 12.070 56.385 12.760 ;
        RECT 59.370 12.070 59.540 12.760 ;
        RECT 60.160 12.070 60.330 12.760 ;
        RECT 60.750 12.070 60.920 12.760 ;
        RECT 61.540 12.070 61.710 12.760 ;
        RECT 64.705 12.070 64.875 12.760 ;
        RECT 65.495 12.070 65.665 12.760 ;
        RECT 66.085 12.070 66.255 12.760 ;
        RECT 66.875 12.070 67.045 12.760 ;
        RECT 70.030 12.070 70.200 12.760 ;
        RECT 70.820 12.070 70.990 12.760 ;
        RECT 71.410 12.070 71.580 12.760 ;
        RECT 72.200 12.070 72.370 12.760 ;
        RECT 75.365 12.070 75.535 12.760 ;
        RECT 76.155 12.070 76.325 12.760 ;
        RECT 76.745 12.070 76.915 12.760 ;
        RECT 77.535 12.070 77.705 12.760 ;
        RECT 80.690 12.070 80.860 12.760 ;
        RECT 81.480 12.070 81.650 12.760 ;
        RECT 82.070 12.070 82.240 12.760 ;
        RECT 82.860 12.070 83.030 12.760 ;
        RECT 86.025 12.070 86.195 12.760 ;
        RECT 86.815 12.070 86.985 12.760 ;
        RECT 87.405 12.070 87.575 12.760 ;
        RECT 88.195 12.070 88.365 12.760 ;
        RECT 91.350 12.070 91.520 12.760 ;
        RECT 92.140 12.070 92.310 12.760 ;
        RECT 92.730 12.070 92.900 12.760 ;
        RECT 93.520 12.070 93.690 12.760 ;
        RECT 96.685 12.070 96.855 12.760 ;
        RECT 97.475 12.070 97.645 12.760 ;
        RECT 98.065 12.070 98.235 12.760 ;
        RECT 98.855 12.070 99.025 12.760 ;
        RECT 102.010 12.070 102.180 12.760 ;
        RECT 102.800 12.070 102.970 12.760 ;
        RECT 103.390 12.070 103.560 12.760 ;
        RECT 104.180 12.070 104.350 12.760 ;
        RECT 107.345 12.070 107.515 12.760 ;
        RECT 108.135 12.070 108.305 12.760 ;
        RECT 108.725 12.070 108.895 12.760 ;
        RECT 109.515 12.070 109.685 12.760 ;
        RECT 112.670 12.070 112.840 12.760 ;
        RECT 113.460 12.070 113.630 12.760 ;
        RECT 114.050 12.070 114.220 12.760 ;
        RECT 114.840 12.070 115.010 12.760 ;
        RECT 118.005 12.070 118.175 12.760 ;
        RECT 118.795 12.070 118.965 12.760 ;
        RECT 119.385 12.070 119.555 12.760 ;
        RECT 120.175 12.070 120.345 12.760 ;
        RECT 124.120 12.070 124.290 12.760 ;
        RECT 124.710 12.070 124.880 12.760 ;
        RECT 125.500 12.070 125.670 12.760 ;
        RECT 16.175 11.910 20.400 11.925 ;
        RECT 14.645 11.705 15.945 11.735 ;
        RECT 12.130 11.500 12.685 11.670 ;
        RECT 12.455 11.260 12.685 11.500 ;
        RECT 13.600 11.470 20.050 11.705 ;
        RECT 12.090 10.430 12.685 11.260 ;
        RECT 14.485 11.285 19.515 11.290 ;
        RECT 20.230 11.285 20.400 11.910 ;
        RECT 14.485 11.120 20.400 11.285 ;
        RECT 14.485 10.620 14.695 11.120 ;
        RECT 16.045 11.115 20.400 11.120 ;
        RECT 16.045 11.105 20.260 11.115 ;
        RECT 16.045 10.620 16.255 11.105 ;
        RECT 17.605 10.620 17.815 11.105 ;
        RECT 19.205 10.620 19.855 11.105 ;
        RECT 2.825 7.745 3.155 9.295 ;
        RECT 4.385 7.745 4.715 9.295 ;
        RECT 5.945 7.745 6.275 9.375 ;
        RECT 8.845 8.305 9.175 9.375 ;
        RECT 10.450 8.475 10.780 9.375 ;
        RECT 11.930 8.660 12.180 9.395 ;
        RECT 13.490 8.660 14.075 9.395 ;
        RECT 11.930 8.490 14.075 8.660 ;
        RECT 15.925 8.665 16.135 9.160 ;
        RECT 17.485 8.665 17.695 9.160 ;
        RECT 19.045 8.665 19.255 9.160 ;
        RECT 20.645 8.665 21.295 9.160 ;
        RECT 15.925 8.490 21.840 8.665 ;
        RECT 7.990 7.745 8.320 8.305 ;
        RECT 2.825 7.415 8.320 7.745 ;
        RECT 3.215 4.805 3.505 7.245 ;
        RECT 6.515 5.215 6.845 7.415 ;
        RECT 7.990 6.955 8.320 7.415 ;
        RECT 8.845 7.975 10.370 8.305 ;
        RECT 7.015 6.220 7.825 6.550 ;
        RECT 7.495 5.555 7.825 6.220 ;
        RECT 8.845 6.155 9.175 7.975 ;
        RECT 10.540 7.805 10.780 8.475 ;
        RECT 13.905 8.340 14.075 8.490 ;
        RECT 13.905 8.310 14.605 8.340 ;
        RECT 11.015 8.140 13.725 8.310 ;
        RECT 13.905 8.075 21.490 8.310 ;
        RECT 13.905 7.960 15.710 8.075 ;
        RECT 10.450 6.155 10.780 7.805 ;
        RECT 11.930 7.790 15.710 7.960 ;
        RECT 21.670 7.860 21.840 8.490 ;
        RECT 16.045 7.855 21.840 7.860 ;
        RECT 11.930 6.135 12.260 7.790 ;
        RECT 13.570 6.135 13.820 7.790 ;
        RECT 16.005 7.685 21.840 7.855 ;
        RECT 16.005 6.445 16.335 7.685 ;
        RECT 17.565 6.445 17.895 7.685 ;
        RECT 19.125 6.445 19.455 7.685 ;
        RECT 20.685 6.445 21.015 7.685 ;
        RECT 31.475 7.280 32.185 11.855 ;
        RECT 32.725 10.275 32.895 11.315 ;
        RECT 33.515 10.275 33.685 11.315 ;
        RECT 34.105 10.275 34.275 11.315 ;
        RECT 34.895 10.275 35.065 11.315 ;
        RECT 38.840 10.275 39.010 11.315 ;
        RECT 39.430 10.275 39.600 11.315 ;
        RECT 40.220 10.275 40.390 11.315 ;
        RECT 38.280 9.890 38.780 10.060 ;
        RECT 39.660 9.890 40.160 10.060 ;
        RECT 32.725 7.720 32.895 8.760 ;
        RECT 33.515 7.720 33.685 8.760 ;
        RECT 34.105 7.720 34.275 8.760 ;
        RECT 38.050 7.720 38.220 8.760 ;
        RECT 38.840 7.720 39.010 8.760 ;
        RECT 39.430 7.720 39.600 8.760 ;
        RECT 40.220 7.720 40.390 8.760 ;
        RECT 40.935 7.260 41.645 11.835 ;
        RECT 42.135 7.265 42.845 11.840 ;
        RECT 43.385 10.275 43.555 11.315 ;
        RECT 44.175 10.275 44.345 11.315 ;
        RECT 44.765 10.275 44.935 11.315 ;
        RECT 45.555 10.275 45.725 11.315 ;
        RECT 43.615 9.890 44.115 10.060 ;
        RECT 44.995 9.890 45.495 10.060 ;
        RECT 43.385 7.720 43.555 8.760 ;
        RECT 44.175 7.720 44.345 8.760 ;
        RECT 44.765 7.720 44.935 8.760 ;
        RECT 45.555 7.720 45.725 8.760 ;
        RECT 46.270 7.260 46.980 11.835 ;
        RECT 47.460 7.265 48.170 11.840 ;
        RECT 48.710 10.275 48.880 11.315 ;
        RECT 49.500 10.275 49.670 11.315 ;
        RECT 50.090 10.275 50.260 11.315 ;
        RECT 50.880 10.275 51.050 11.315 ;
        RECT 48.940 9.890 49.440 10.060 ;
        RECT 50.320 9.890 50.820 10.060 ;
        RECT 48.710 7.720 48.880 8.760 ;
        RECT 49.500 7.720 49.670 8.760 ;
        RECT 50.090 7.720 50.260 8.760 ;
        RECT 50.880 7.720 51.050 8.760 ;
        RECT 51.595 7.260 52.305 11.835 ;
        RECT 52.795 7.265 53.505 11.840 ;
        RECT 54.045 10.275 54.215 11.315 ;
        RECT 54.835 10.275 55.005 11.315 ;
        RECT 55.425 10.275 55.595 11.315 ;
        RECT 56.215 10.275 56.385 11.315 ;
        RECT 54.275 9.890 54.775 10.060 ;
        RECT 55.655 9.890 56.155 10.060 ;
        RECT 54.045 7.720 54.215 8.760 ;
        RECT 54.835 7.720 55.005 8.760 ;
        RECT 55.425 7.720 55.595 8.760 ;
        RECT 56.215 7.720 56.385 8.760 ;
        RECT 56.930 7.260 57.640 11.835 ;
        RECT 58.120 7.265 58.830 11.840 ;
        RECT 59.370 10.275 59.540 11.315 ;
        RECT 60.160 10.275 60.330 11.315 ;
        RECT 60.750 10.275 60.920 11.315 ;
        RECT 61.540 10.275 61.710 11.315 ;
        RECT 59.600 9.890 60.100 10.060 ;
        RECT 60.980 9.890 61.480 10.060 ;
        RECT 59.370 7.720 59.540 8.760 ;
        RECT 60.160 7.720 60.330 8.760 ;
        RECT 60.750 7.720 60.920 8.760 ;
        RECT 61.540 7.720 61.710 8.760 ;
        RECT 62.255 7.260 62.965 11.835 ;
        RECT 63.455 7.265 64.165 11.840 ;
        RECT 64.705 10.275 64.875 11.315 ;
        RECT 65.495 10.275 65.665 11.315 ;
        RECT 66.085 10.275 66.255 11.315 ;
        RECT 66.875 10.275 67.045 11.315 ;
        RECT 64.935 9.890 65.435 10.060 ;
        RECT 66.315 9.890 66.815 10.060 ;
        RECT 64.705 7.720 64.875 8.760 ;
        RECT 65.495 7.720 65.665 8.760 ;
        RECT 66.085 7.720 66.255 8.760 ;
        RECT 66.875 7.720 67.045 8.760 ;
        RECT 67.590 7.260 68.300 11.835 ;
        RECT 68.780 7.265 69.490 11.840 ;
        RECT 70.030 10.275 70.200 11.315 ;
        RECT 70.820 10.275 70.990 11.315 ;
        RECT 71.410 10.275 71.580 11.315 ;
        RECT 72.200 10.275 72.370 11.315 ;
        RECT 70.260 9.890 70.760 10.060 ;
        RECT 71.640 9.890 72.140 10.060 ;
        RECT 70.030 7.720 70.200 8.760 ;
        RECT 70.820 7.720 70.990 8.760 ;
        RECT 71.410 7.720 71.580 8.760 ;
        RECT 72.200 7.720 72.370 8.760 ;
        RECT 72.915 7.260 73.625 11.835 ;
        RECT 74.115 7.265 74.825 11.840 ;
        RECT 75.365 10.275 75.535 11.315 ;
        RECT 76.155 10.275 76.325 11.315 ;
        RECT 76.745 10.275 76.915 11.315 ;
        RECT 77.535 10.275 77.705 11.315 ;
        RECT 75.595 9.890 76.095 10.060 ;
        RECT 76.975 9.890 77.475 10.060 ;
        RECT 75.365 7.720 75.535 8.760 ;
        RECT 76.155 7.720 76.325 8.760 ;
        RECT 76.745 7.720 76.915 8.760 ;
        RECT 77.535 7.720 77.705 8.760 ;
        RECT 78.250 7.260 78.960 11.835 ;
        RECT 79.440 7.265 80.150 11.840 ;
        RECT 80.690 10.275 80.860 11.315 ;
        RECT 81.480 10.275 81.650 11.315 ;
        RECT 82.070 10.275 82.240 11.315 ;
        RECT 82.860 10.275 83.030 11.315 ;
        RECT 80.920 9.890 81.420 10.060 ;
        RECT 82.300 9.890 82.800 10.060 ;
        RECT 80.690 7.720 80.860 8.760 ;
        RECT 81.480 7.720 81.650 8.760 ;
        RECT 82.070 7.720 82.240 8.760 ;
        RECT 82.860 7.720 83.030 8.760 ;
        RECT 83.575 7.260 84.285 11.835 ;
        RECT 84.775 7.265 85.485 11.840 ;
        RECT 86.025 10.275 86.195 11.315 ;
        RECT 86.815 10.275 86.985 11.315 ;
        RECT 87.405 10.275 87.575 11.315 ;
        RECT 88.195 10.275 88.365 11.315 ;
        RECT 86.255 9.890 86.755 10.060 ;
        RECT 87.635 9.890 88.135 10.060 ;
        RECT 86.025 7.720 86.195 8.760 ;
        RECT 86.815 7.720 86.985 8.760 ;
        RECT 87.405 7.720 87.575 8.760 ;
        RECT 88.195 7.720 88.365 8.760 ;
        RECT 88.910 7.260 89.620 11.835 ;
        RECT 90.100 7.265 90.810 11.840 ;
        RECT 91.350 10.275 91.520 11.315 ;
        RECT 92.140 10.275 92.310 11.315 ;
        RECT 92.730 10.275 92.900 11.315 ;
        RECT 93.520 10.275 93.690 11.315 ;
        RECT 91.580 9.890 92.080 10.060 ;
        RECT 92.960 9.890 93.460 10.060 ;
        RECT 91.350 7.720 91.520 8.760 ;
        RECT 92.140 7.720 92.310 8.760 ;
        RECT 92.730 7.720 92.900 8.760 ;
        RECT 93.520 7.720 93.690 8.760 ;
        RECT 94.235 7.260 94.945 11.835 ;
        RECT 95.435 7.265 96.145 11.840 ;
        RECT 96.685 10.275 96.855 11.315 ;
        RECT 97.475 10.275 97.645 11.315 ;
        RECT 98.065 10.275 98.235 11.315 ;
        RECT 98.855 10.275 99.025 11.315 ;
        RECT 96.915 9.890 97.415 10.060 ;
        RECT 98.295 9.890 98.795 10.060 ;
        RECT 96.685 7.720 96.855 8.760 ;
        RECT 97.475 7.720 97.645 8.760 ;
        RECT 98.065 7.720 98.235 8.760 ;
        RECT 98.855 7.720 99.025 8.760 ;
        RECT 99.570 7.260 100.280 11.835 ;
        RECT 100.760 7.265 101.470 11.840 ;
        RECT 102.010 10.275 102.180 11.315 ;
        RECT 102.800 10.275 102.970 11.315 ;
        RECT 103.390 10.275 103.560 11.315 ;
        RECT 104.180 10.275 104.350 11.315 ;
        RECT 102.240 9.890 102.740 10.060 ;
        RECT 103.620 9.890 104.120 10.060 ;
        RECT 102.010 7.720 102.180 8.760 ;
        RECT 102.800 7.720 102.970 8.760 ;
        RECT 103.390 7.720 103.560 8.760 ;
        RECT 104.180 7.720 104.350 8.760 ;
        RECT 104.895 7.260 105.605 11.835 ;
        RECT 106.095 7.265 106.805 11.840 ;
        RECT 107.345 10.275 107.515 11.315 ;
        RECT 108.135 10.275 108.305 11.315 ;
        RECT 108.725 10.275 108.895 11.315 ;
        RECT 109.515 10.275 109.685 11.315 ;
        RECT 107.575 9.890 108.075 10.060 ;
        RECT 108.955 9.890 109.455 10.060 ;
        RECT 107.345 7.720 107.515 8.760 ;
        RECT 108.135 7.720 108.305 8.760 ;
        RECT 108.725 7.720 108.895 8.760 ;
        RECT 109.515 7.720 109.685 8.760 ;
        RECT 110.230 7.260 110.940 11.835 ;
        RECT 111.420 7.265 112.130 11.840 ;
        RECT 112.670 10.275 112.840 11.315 ;
        RECT 113.460 10.275 113.630 11.315 ;
        RECT 114.050 10.275 114.220 11.315 ;
        RECT 114.840 10.275 115.010 11.315 ;
        RECT 112.900 9.890 113.400 10.060 ;
        RECT 114.280 9.890 114.780 10.060 ;
        RECT 112.670 7.720 112.840 8.760 ;
        RECT 113.460 7.720 113.630 8.760 ;
        RECT 114.050 7.720 114.220 8.760 ;
        RECT 114.840 7.720 115.010 8.760 ;
        RECT 115.555 7.260 116.265 11.835 ;
        RECT 116.755 7.265 117.465 11.840 ;
        RECT 118.005 10.275 118.175 11.315 ;
        RECT 118.795 10.275 118.965 11.315 ;
        RECT 119.385 10.275 119.555 11.315 ;
        RECT 120.175 10.275 120.345 11.315 ;
        RECT 124.120 10.275 124.290 11.315 ;
        RECT 124.710 10.275 124.880 11.315 ;
        RECT 125.500 10.275 125.670 11.315 ;
        RECT 118.235 9.890 118.735 10.060 ;
        RECT 119.615 9.890 120.115 10.060 ;
        RECT 118.005 7.720 118.175 8.760 ;
        RECT 118.795 7.720 118.965 8.760 ;
        RECT 119.385 7.720 119.555 8.760 ;
        RECT 123.330 7.720 123.500 8.760 ;
        RECT 124.120 7.720 124.290 8.760 ;
        RECT 124.710 7.720 124.880 8.760 ;
        RECT 125.500 7.720 125.670 8.760 ;
        RECT 126.215 7.280 126.925 11.855 ;
        RECT 32.725 6.275 32.895 6.965 ;
        RECT 33.515 6.275 33.685 6.965 ;
        RECT 34.105 6.275 34.275 6.965 ;
        RECT 38.050 6.275 38.220 6.965 ;
        RECT 38.840 6.275 39.010 6.965 ;
        RECT 39.430 6.275 39.600 6.965 ;
        RECT 40.220 6.275 40.390 6.965 ;
        RECT 43.385 6.275 43.555 6.965 ;
        RECT 44.175 6.275 44.345 6.965 ;
        RECT 44.765 6.275 44.935 6.965 ;
        RECT 45.555 6.275 45.725 6.965 ;
        RECT 48.710 6.275 48.880 6.965 ;
        RECT 49.500 6.275 49.670 6.965 ;
        RECT 50.090 6.275 50.260 6.965 ;
        RECT 50.880 6.275 51.050 6.965 ;
        RECT 54.045 6.275 54.215 6.965 ;
        RECT 54.835 6.275 55.005 6.965 ;
        RECT 55.425 6.275 55.595 6.965 ;
        RECT 56.215 6.275 56.385 6.965 ;
        RECT 59.370 6.275 59.540 6.965 ;
        RECT 60.160 6.275 60.330 6.965 ;
        RECT 60.750 6.275 60.920 6.965 ;
        RECT 61.540 6.275 61.710 6.965 ;
        RECT 64.705 6.275 64.875 6.965 ;
        RECT 65.495 6.275 65.665 6.965 ;
        RECT 66.085 6.275 66.255 6.965 ;
        RECT 66.875 6.275 67.045 6.965 ;
        RECT 70.030 6.275 70.200 6.965 ;
        RECT 70.820 6.275 70.990 6.965 ;
        RECT 71.410 6.275 71.580 6.965 ;
        RECT 72.200 6.275 72.370 6.965 ;
        RECT 75.365 6.275 75.535 6.965 ;
        RECT 76.155 6.275 76.325 6.965 ;
        RECT 76.745 6.275 76.915 6.965 ;
        RECT 77.535 6.275 77.705 6.965 ;
        RECT 80.690 6.275 80.860 6.965 ;
        RECT 81.480 6.275 81.650 6.965 ;
        RECT 82.070 6.275 82.240 6.965 ;
        RECT 82.860 6.275 83.030 6.965 ;
        RECT 86.025 6.275 86.195 6.965 ;
        RECT 86.815 6.275 86.985 6.965 ;
        RECT 87.405 6.275 87.575 6.965 ;
        RECT 88.195 6.275 88.365 6.965 ;
        RECT 91.350 6.275 91.520 6.965 ;
        RECT 92.140 6.275 92.310 6.965 ;
        RECT 92.730 6.275 92.900 6.965 ;
        RECT 93.520 6.275 93.690 6.965 ;
        RECT 96.685 6.275 96.855 6.965 ;
        RECT 97.475 6.275 97.645 6.965 ;
        RECT 98.065 6.275 98.235 6.965 ;
        RECT 98.855 6.275 99.025 6.965 ;
        RECT 102.010 6.275 102.180 6.965 ;
        RECT 102.800 6.275 102.970 6.965 ;
        RECT 103.390 6.275 103.560 6.965 ;
        RECT 104.180 6.275 104.350 6.965 ;
        RECT 107.345 6.275 107.515 6.965 ;
        RECT 108.135 6.275 108.305 6.965 ;
        RECT 108.725 6.275 108.895 6.965 ;
        RECT 109.515 6.275 109.685 6.965 ;
        RECT 112.670 6.275 112.840 6.965 ;
        RECT 113.460 6.275 113.630 6.965 ;
        RECT 114.050 6.275 114.220 6.965 ;
        RECT 114.840 6.275 115.010 6.965 ;
        RECT 118.005 6.275 118.175 6.965 ;
        RECT 118.795 6.275 118.965 6.965 ;
        RECT 119.385 6.275 119.555 6.965 ;
        RECT 123.330 6.275 123.500 6.965 ;
        RECT 124.120 6.275 124.290 6.965 ;
        RECT 124.710 6.275 124.880 6.965 ;
        RECT 125.500 6.275 125.670 6.965 ;
        RECT 6.515 4.885 7.325 5.215 ;
        RECT 3.215 4.515 3.595 4.805 ;
        RECT 3.305 3.745 3.595 4.515 ;
        RECT 4.205 4.225 4.515 4.655 ;
        RECT 6.995 4.545 7.325 4.885 ;
        RECT 7.495 5.145 8.165 5.555 ;
        RECT 7.495 4.225 7.825 5.145 ;
        RECT 4.205 3.915 6.120 4.225 ;
        RECT 4.810 3.895 6.120 3.915 ;
        RECT 6.290 3.895 9.740 4.225 ;
        RECT 3.305 3.495 4.640 3.745 ;
        RECT 3.305 2.485 3.595 3.495 ;
        RECT 4.810 3.325 5.140 3.895 ;
        RECT 4.205 2.995 5.140 3.325 ;
        RECT 4.205 2.485 4.515 2.995 ;
        RECT 6.290 2.345 6.620 3.895 ;
        RECT 7.850 2.345 8.180 3.895 ;
        RECT 9.410 2.265 9.740 3.895 ;
        RECT 11.015 3.300 11.960 3.630 ;
        RECT 12.130 3.530 12.380 5.505 ;
        RECT 14.565 3.955 14.895 5.195 ;
        RECT 16.125 3.955 16.455 5.195 ;
        RECT 17.685 3.955 18.015 5.195 ;
        RECT 19.245 3.955 19.575 5.195 ;
        RECT 32.725 4.535 32.895 5.225 ;
        RECT 33.515 4.535 33.685 5.225 ;
        RECT 34.105 4.535 34.275 5.225 ;
        RECT 34.895 4.535 35.065 5.225 ;
        RECT 38.050 4.535 38.220 5.225 ;
        RECT 38.840 4.535 39.010 5.225 ;
        RECT 39.430 4.535 39.600 5.225 ;
        RECT 40.220 4.535 40.390 5.225 ;
        RECT 43.385 4.535 43.555 5.225 ;
        RECT 44.175 4.535 44.345 5.225 ;
        RECT 44.765 4.535 44.935 5.225 ;
        RECT 45.555 4.535 45.725 5.225 ;
        RECT 48.710 4.535 48.880 5.225 ;
        RECT 49.500 4.535 49.670 5.225 ;
        RECT 50.090 4.535 50.260 5.225 ;
        RECT 50.880 4.535 51.050 5.225 ;
        RECT 54.045 4.535 54.215 5.225 ;
        RECT 54.835 4.535 55.005 5.225 ;
        RECT 55.425 4.535 55.595 5.225 ;
        RECT 56.215 4.535 56.385 5.225 ;
        RECT 59.370 4.535 59.540 5.225 ;
        RECT 60.160 4.535 60.330 5.225 ;
        RECT 60.750 4.535 60.920 5.225 ;
        RECT 61.540 4.535 61.710 5.225 ;
        RECT 64.705 4.535 64.875 5.225 ;
        RECT 65.495 4.535 65.665 5.225 ;
        RECT 66.085 4.535 66.255 5.225 ;
        RECT 66.875 4.535 67.045 5.225 ;
        RECT 70.030 4.535 70.200 5.225 ;
        RECT 70.820 4.535 70.990 5.225 ;
        RECT 71.410 4.535 71.580 5.225 ;
        RECT 72.200 4.535 72.370 5.225 ;
        RECT 75.365 4.535 75.535 5.225 ;
        RECT 76.155 4.535 76.325 5.225 ;
        RECT 76.745 4.535 76.915 5.225 ;
        RECT 77.535 4.535 77.705 5.225 ;
        RECT 80.690 4.535 80.860 5.225 ;
        RECT 81.480 4.535 81.650 5.225 ;
        RECT 82.070 4.535 82.240 5.225 ;
        RECT 82.860 4.535 83.030 5.225 ;
        RECT 86.025 4.535 86.195 5.225 ;
        RECT 86.815 4.535 86.985 5.225 ;
        RECT 87.405 4.535 87.575 5.225 ;
        RECT 88.195 4.535 88.365 5.225 ;
        RECT 91.350 4.535 91.520 5.225 ;
        RECT 92.140 4.535 92.310 5.225 ;
        RECT 92.730 4.535 92.900 5.225 ;
        RECT 93.520 4.535 93.690 5.225 ;
        RECT 96.685 4.535 96.855 5.225 ;
        RECT 97.475 4.535 97.645 5.225 ;
        RECT 98.065 4.535 98.235 5.225 ;
        RECT 98.855 4.535 99.025 5.225 ;
        RECT 102.010 4.535 102.180 5.225 ;
        RECT 102.800 4.535 102.970 5.225 ;
        RECT 103.390 4.535 103.560 5.225 ;
        RECT 104.180 4.535 104.350 5.225 ;
        RECT 107.345 4.535 107.515 5.225 ;
        RECT 108.135 4.535 108.305 5.225 ;
        RECT 108.725 4.535 108.895 5.225 ;
        RECT 109.515 4.535 109.685 5.225 ;
        RECT 112.670 4.535 112.840 5.225 ;
        RECT 113.460 4.535 113.630 5.225 ;
        RECT 114.050 4.535 114.220 5.225 ;
        RECT 114.840 4.535 115.010 5.225 ;
        RECT 118.005 4.535 118.175 5.225 ;
        RECT 118.795 4.535 118.965 5.225 ;
        RECT 119.385 4.535 119.555 5.225 ;
        RECT 120.175 4.535 120.345 5.225 ;
        RECT 123.330 4.535 123.500 5.225 ;
        RECT 124.120 4.535 124.290 5.225 ;
        RECT 124.710 4.535 124.880 5.225 ;
        RECT 125.500 4.535 125.670 5.225 ;
        RECT 14.565 3.785 20.400 3.955 ;
        RECT 16.175 3.770 20.400 3.785 ;
        RECT 14.645 3.565 15.945 3.595 ;
        RECT 12.130 3.360 12.685 3.530 ;
        RECT 12.455 3.120 12.685 3.360 ;
        RECT 13.600 3.330 20.050 3.565 ;
        RECT 12.090 2.290 12.685 3.120 ;
        RECT 14.485 3.145 19.515 3.150 ;
        RECT 20.230 3.145 20.400 3.770 ;
        RECT 14.485 2.980 20.400 3.145 ;
        RECT 14.485 2.480 14.695 2.980 ;
        RECT 16.045 2.975 20.400 2.980 ;
        RECT 16.045 2.965 20.260 2.975 ;
        RECT 16.045 2.480 16.255 2.965 ;
        RECT 17.605 2.480 17.815 2.965 ;
        RECT 19.205 2.480 19.855 2.965 ;
        RECT 31.475 2.030 32.185 4.320 ;
        RECT 32.725 2.740 32.895 3.780 ;
        RECT 33.515 2.740 33.685 3.780 ;
        RECT 34.105 2.740 34.275 3.780 ;
        RECT 34.895 2.740 35.065 3.780 ;
        RECT 35.610 2.030 36.320 4.320 ;
        RECT 36.800 2.015 37.510 4.305 ;
        RECT 38.050 2.740 38.220 3.780 ;
        RECT 38.840 2.740 39.010 3.780 ;
        RECT 39.430 2.740 39.600 3.780 ;
        RECT 40.220 2.740 40.390 3.780 ;
        RECT 40.935 2.010 41.645 4.300 ;
        RECT 42.135 2.015 42.845 4.305 ;
        RECT 43.385 2.740 43.555 3.780 ;
        RECT 44.175 2.740 44.345 3.780 ;
        RECT 44.765 2.740 44.935 3.780 ;
        RECT 45.555 2.740 45.725 3.780 ;
        RECT 46.270 2.010 46.980 4.300 ;
        RECT 47.460 2.015 48.170 4.305 ;
        RECT 48.710 2.740 48.880 3.780 ;
        RECT 49.500 2.740 49.670 3.780 ;
        RECT 50.090 2.740 50.260 3.780 ;
        RECT 50.880 2.740 51.050 3.780 ;
        RECT 51.595 2.010 52.305 4.300 ;
        RECT 52.795 2.015 53.505 4.305 ;
        RECT 54.045 2.740 54.215 3.780 ;
        RECT 54.835 2.740 55.005 3.780 ;
        RECT 55.425 2.740 55.595 3.780 ;
        RECT 56.215 2.740 56.385 3.780 ;
        RECT 56.930 2.010 57.640 4.300 ;
        RECT 58.120 2.015 58.830 4.305 ;
        RECT 59.370 2.740 59.540 3.780 ;
        RECT 60.160 2.740 60.330 3.780 ;
        RECT 60.750 2.740 60.920 3.780 ;
        RECT 61.540 2.740 61.710 3.780 ;
        RECT 62.255 2.010 62.965 4.300 ;
        RECT 63.455 2.015 64.165 4.305 ;
        RECT 64.705 2.740 64.875 3.780 ;
        RECT 65.495 2.740 65.665 3.780 ;
        RECT 66.085 2.740 66.255 3.780 ;
        RECT 66.875 2.740 67.045 3.780 ;
        RECT 67.590 2.010 68.300 4.300 ;
        RECT 68.780 2.015 69.490 4.305 ;
        RECT 70.030 2.740 70.200 3.780 ;
        RECT 70.820 2.740 70.990 3.780 ;
        RECT 71.410 2.740 71.580 3.780 ;
        RECT 72.200 2.740 72.370 3.780 ;
        RECT 72.915 2.010 73.625 4.300 ;
        RECT 74.115 2.015 74.825 4.305 ;
        RECT 75.365 2.740 75.535 3.780 ;
        RECT 76.155 2.740 76.325 3.780 ;
        RECT 76.745 2.740 76.915 3.780 ;
        RECT 77.535 2.740 77.705 3.780 ;
        RECT 78.250 2.010 78.960 4.300 ;
        RECT 79.440 2.015 80.150 4.305 ;
        RECT 80.690 2.740 80.860 3.780 ;
        RECT 81.480 2.740 81.650 3.780 ;
        RECT 82.070 2.740 82.240 3.780 ;
        RECT 82.860 2.740 83.030 3.780 ;
        RECT 83.575 2.010 84.285 4.300 ;
        RECT 84.775 2.015 85.485 4.305 ;
        RECT 86.025 2.740 86.195 3.780 ;
        RECT 86.815 2.740 86.985 3.780 ;
        RECT 87.405 2.740 87.575 3.780 ;
        RECT 88.195 2.740 88.365 3.780 ;
        RECT 88.910 2.010 89.620 4.300 ;
        RECT 90.100 2.015 90.810 4.305 ;
        RECT 91.350 2.740 91.520 3.780 ;
        RECT 92.140 2.740 92.310 3.780 ;
        RECT 92.730 2.740 92.900 3.780 ;
        RECT 93.520 2.740 93.690 3.780 ;
        RECT 94.235 2.010 94.945 4.300 ;
        RECT 95.435 2.015 96.145 4.305 ;
        RECT 96.685 2.740 96.855 3.780 ;
        RECT 97.475 2.740 97.645 3.780 ;
        RECT 98.065 2.740 98.235 3.780 ;
        RECT 98.855 2.740 99.025 3.780 ;
        RECT 99.570 2.010 100.280 4.300 ;
        RECT 100.760 2.015 101.470 4.305 ;
        RECT 102.010 2.740 102.180 3.780 ;
        RECT 102.800 2.740 102.970 3.780 ;
        RECT 103.390 2.740 103.560 3.780 ;
        RECT 104.180 2.740 104.350 3.780 ;
        RECT 104.895 2.010 105.605 4.300 ;
        RECT 106.095 2.015 106.805 4.305 ;
        RECT 107.345 2.740 107.515 3.780 ;
        RECT 108.135 2.740 108.305 3.780 ;
        RECT 108.725 2.740 108.895 3.780 ;
        RECT 109.515 2.740 109.685 3.780 ;
        RECT 110.230 2.010 110.940 4.300 ;
        RECT 111.420 2.015 112.130 4.305 ;
        RECT 112.670 2.740 112.840 3.780 ;
        RECT 113.460 2.740 113.630 3.780 ;
        RECT 114.050 2.740 114.220 3.780 ;
        RECT 114.840 2.740 115.010 3.780 ;
        RECT 115.555 2.010 116.265 4.300 ;
        RECT 116.755 2.015 117.465 4.305 ;
        RECT 118.005 2.740 118.175 3.780 ;
        RECT 118.795 2.740 118.965 3.780 ;
        RECT 119.385 2.740 119.555 3.780 ;
        RECT 120.175 2.740 120.345 3.780 ;
        RECT 120.890 2.010 121.600 4.300 ;
        RECT 122.080 2.030 122.790 4.320 ;
        RECT 123.330 2.740 123.500 3.780 ;
        RECT 124.120 2.740 124.290 3.780 ;
        RECT 124.710 2.740 124.880 3.780 ;
        RECT 125.500 2.740 125.670 3.780 ;
        RECT 126.215 2.030 126.925 4.320 ;
      LAYER met1 ;
        RECT 32.635 77.705 35.185 77.970 ;
        RECT 32.635 77.500 32.970 77.705 ;
        RECT 31.470 77.380 32.970 77.500 ;
        RECT 31.420 77.185 32.970 77.380 ;
        RECT 34.850 77.460 35.185 77.705 ;
        RECT 38.515 77.690 39.930 77.930 ;
        RECT 34.850 77.380 36.270 77.460 ;
        RECT 38.515 77.425 38.755 77.690 ;
        RECT 34.850 77.185 36.375 77.380 ;
        RECT 36.845 77.365 38.755 77.425 ;
        RECT 31.420 77.165 31.820 77.185 ;
        RECT 31.420 75.095 31.775 77.165 ;
        RECT 32.695 75.320 32.925 76.555 ;
        RECT 33.485 75.320 33.715 76.555 ;
        RECT 34.075 75.320 34.305 76.555 ;
        RECT 32.680 75.000 32.940 75.320 ;
        RECT 33.470 75.000 33.730 75.320 ;
        RECT 34.060 75.000 34.320 75.320 ;
        RECT 34.865 75.245 35.095 76.555 ;
        RECT 35.705 75.245 35.875 77.185 ;
        RECT 34.865 75.075 35.875 75.245 ;
        RECT 36.020 75.095 36.375 77.185 ;
        RECT 36.745 77.185 38.755 77.365 ;
        RECT 39.690 77.460 39.930 77.690 ;
        RECT 43.845 77.685 45.255 77.925 ;
        RECT 39.690 77.360 41.595 77.460 ;
        RECT 43.845 77.425 44.085 77.685 ;
        RECT 42.180 77.365 44.085 77.425 ;
        RECT 39.690 77.220 41.700 77.360 ;
        RECT 41.030 77.185 41.700 77.220 ;
        RECT 36.745 75.080 37.100 77.185 ;
        RECT 38.020 75.320 38.250 76.555 ;
        RECT 38.810 75.320 39.040 76.555 ;
        RECT 39.400 75.320 39.630 76.555 ;
        RECT 32.695 74.110 32.925 75.000 ;
        RECT 33.485 74.110 33.715 75.000 ;
        RECT 34.075 74.110 34.305 75.000 ;
        RECT 34.865 74.110 35.095 75.075 ;
        RECT 38.005 75.000 38.265 75.320 ;
        RECT 38.795 75.000 39.055 75.320 ;
        RECT 39.385 75.000 39.645 75.320 ;
        RECT 40.190 75.245 40.420 76.555 ;
        RECT 41.030 75.245 41.200 77.185 ;
        RECT 40.190 75.075 41.200 75.245 ;
        RECT 41.345 75.075 41.700 77.185 ;
        RECT 42.080 77.185 44.085 77.365 ;
        RECT 45.015 77.460 45.255 77.685 ;
        RECT 49.175 77.690 50.590 77.930 ;
        RECT 45.015 77.360 46.930 77.460 ;
        RECT 49.175 77.425 49.415 77.690 ;
        RECT 47.505 77.365 49.415 77.425 ;
        RECT 45.015 77.220 47.035 77.360 ;
        RECT 46.365 77.185 47.035 77.220 ;
        RECT 42.080 75.080 42.435 77.185 ;
        RECT 43.355 75.320 43.585 76.555 ;
        RECT 44.145 75.320 44.375 76.555 ;
        RECT 44.735 75.320 44.965 76.555 ;
        RECT 38.020 74.110 38.250 75.000 ;
        RECT 38.810 74.110 39.040 75.000 ;
        RECT 39.400 74.110 39.630 75.000 ;
        RECT 40.190 74.110 40.420 75.075 ;
        RECT 43.340 75.000 43.600 75.320 ;
        RECT 44.130 75.000 44.390 75.320 ;
        RECT 44.720 75.000 44.980 75.320 ;
        RECT 45.525 75.245 45.755 76.555 ;
        RECT 46.365 75.245 46.535 77.185 ;
        RECT 45.525 75.075 46.535 75.245 ;
        RECT 46.680 75.075 47.035 77.185 ;
        RECT 47.405 77.185 49.415 77.365 ;
        RECT 50.350 77.460 50.590 77.690 ;
        RECT 54.505 77.685 55.915 77.925 ;
        RECT 50.350 77.360 52.255 77.460 ;
        RECT 54.505 77.425 54.745 77.685 ;
        RECT 52.840 77.365 54.745 77.425 ;
        RECT 50.350 77.220 52.360 77.360 ;
        RECT 51.690 77.185 52.360 77.220 ;
        RECT 47.405 75.080 47.760 77.185 ;
        RECT 48.680 75.320 48.910 76.555 ;
        RECT 49.470 75.320 49.700 76.555 ;
        RECT 50.060 75.320 50.290 76.555 ;
        RECT 43.355 74.110 43.585 75.000 ;
        RECT 44.145 74.110 44.375 75.000 ;
        RECT 44.735 74.110 44.965 75.000 ;
        RECT 45.525 74.110 45.755 75.075 ;
        RECT 48.665 75.000 48.925 75.320 ;
        RECT 49.455 75.000 49.715 75.320 ;
        RECT 50.045 75.000 50.305 75.320 ;
        RECT 50.850 75.245 51.080 76.555 ;
        RECT 51.690 75.245 51.860 77.185 ;
        RECT 50.850 75.075 51.860 75.245 ;
        RECT 52.005 75.075 52.360 77.185 ;
        RECT 52.740 77.185 54.745 77.365 ;
        RECT 55.675 77.460 55.915 77.685 ;
        RECT 59.835 77.690 61.250 77.930 ;
        RECT 55.675 77.360 57.590 77.460 ;
        RECT 59.835 77.425 60.075 77.690 ;
        RECT 58.165 77.365 60.075 77.425 ;
        RECT 55.675 77.220 57.695 77.360 ;
        RECT 57.025 77.185 57.695 77.220 ;
        RECT 52.740 75.080 53.095 77.185 ;
        RECT 54.015 75.320 54.245 76.555 ;
        RECT 54.805 75.320 55.035 76.555 ;
        RECT 55.395 75.320 55.625 76.555 ;
        RECT 48.680 74.110 48.910 75.000 ;
        RECT 49.470 74.110 49.700 75.000 ;
        RECT 50.060 74.110 50.290 75.000 ;
        RECT 50.850 74.110 51.080 75.075 ;
        RECT 54.000 75.000 54.260 75.320 ;
        RECT 54.790 75.000 55.050 75.320 ;
        RECT 55.380 75.000 55.640 75.320 ;
        RECT 56.185 75.245 56.415 76.555 ;
        RECT 57.025 75.245 57.195 77.185 ;
        RECT 56.185 75.075 57.195 75.245 ;
        RECT 57.340 75.075 57.695 77.185 ;
        RECT 58.065 77.185 60.075 77.365 ;
        RECT 61.010 77.460 61.250 77.690 ;
        RECT 65.165 77.685 66.575 77.925 ;
        RECT 61.010 77.360 62.915 77.460 ;
        RECT 65.165 77.425 65.405 77.685 ;
        RECT 63.500 77.365 65.405 77.425 ;
        RECT 61.010 77.220 63.020 77.360 ;
        RECT 62.350 77.185 63.020 77.220 ;
        RECT 58.065 75.080 58.420 77.185 ;
        RECT 59.340 75.320 59.570 76.555 ;
        RECT 60.130 75.320 60.360 76.555 ;
        RECT 60.720 75.320 60.950 76.555 ;
        RECT 54.015 74.110 54.245 75.000 ;
        RECT 54.805 74.110 55.035 75.000 ;
        RECT 55.395 74.110 55.625 75.000 ;
        RECT 56.185 74.110 56.415 75.075 ;
        RECT 59.325 75.000 59.585 75.320 ;
        RECT 60.115 75.000 60.375 75.320 ;
        RECT 60.705 75.000 60.965 75.320 ;
        RECT 61.510 75.245 61.740 76.555 ;
        RECT 62.350 75.245 62.520 77.185 ;
        RECT 61.510 75.075 62.520 75.245 ;
        RECT 62.665 75.075 63.020 77.185 ;
        RECT 63.400 77.185 65.405 77.365 ;
        RECT 66.335 77.460 66.575 77.685 ;
        RECT 70.495 77.690 71.910 77.930 ;
        RECT 66.335 77.360 68.250 77.460 ;
        RECT 70.495 77.425 70.735 77.690 ;
        RECT 68.825 77.365 70.735 77.425 ;
        RECT 66.335 77.220 68.355 77.360 ;
        RECT 67.685 77.185 68.355 77.220 ;
        RECT 63.400 75.080 63.755 77.185 ;
        RECT 64.675 75.320 64.905 76.555 ;
        RECT 65.465 75.320 65.695 76.555 ;
        RECT 66.055 75.320 66.285 76.555 ;
        RECT 59.340 74.110 59.570 75.000 ;
        RECT 60.130 74.110 60.360 75.000 ;
        RECT 60.720 74.110 60.950 75.000 ;
        RECT 61.510 74.110 61.740 75.075 ;
        RECT 64.660 75.000 64.920 75.320 ;
        RECT 65.450 75.000 65.710 75.320 ;
        RECT 66.040 75.000 66.300 75.320 ;
        RECT 66.845 75.245 67.075 76.555 ;
        RECT 67.685 75.245 67.855 77.185 ;
        RECT 66.845 75.075 67.855 75.245 ;
        RECT 68.000 75.075 68.355 77.185 ;
        RECT 68.725 77.185 70.735 77.365 ;
        RECT 71.670 77.460 71.910 77.690 ;
        RECT 75.825 77.685 77.235 77.925 ;
        RECT 71.670 77.360 73.575 77.460 ;
        RECT 75.825 77.425 76.065 77.685 ;
        RECT 74.160 77.365 76.065 77.425 ;
        RECT 71.670 77.220 73.680 77.360 ;
        RECT 73.010 77.185 73.680 77.220 ;
        RECT 68.725 75.080 69.080 77.185 ;
        RECT 70.000 75.320 70.230 76.555 ;
        RECT 70.790 75.320 71.020 76.555 ;
        RECT 71.380 75.320 71.610 76.555 ;
        RECT 64.675 74.110 64.905 75.000 ;
        RECT 65.465 74.110 65.695 75.000 ;
        RECT 66.055 74.110 66.285 75.000 ;
        RECT 66.845 74.110 67.075 75.075 ;
        RECT 69.985 75.000 70.245 75.320 ;
        RECT 70.775 75.000 71.035 75.320 ;
        RECT 71.365 75.000 71.625 75.320 ;
        RECT 72.170 75.245 72.400 76.555 ;
        RECT 73.010 75.245 73.180 77.185 ;
        RECT 72.170 75.075 73.180 75.245 ;
        RECT 73.325 75.075 73.680 77.185 ;
        RECT 74.060 77.185 76.065 77.365 ;
        RECT 76.995 77.460 77.235 77.685 ;
        RECT 81.155 77.690 82.570 77.930 ;
        RECT 76.995 77.360 78.910 77.460 ;
        RECT 81.155 77.425 81.395 77.690 ;
        RECT 79.485 77.365 81.395 77.425 ;
        RECT 76.995 77.220 79.015 77.360 ;
        RECT 78.345 77.185 79.015 77.220 ;
        RECT 74.060 75.080 74.415 77.185 ;
        RECT 75.335 75.320 75.565 76.555 ;
        RECT 76.125 75.320 76.355 76.555 ;
        RECT 76.715 75.320 76.945 76.555 ;
        RECT 70.000 74.110 70.230 75.000 ;
        RECT 70.790 74.110 71.020 75.000 ;
        RECT 71.380 74.110 71.610 75.000 ;
        RECT 72.170 74.110 72.400 75.075 ;
        RECT 75.320 75.000 75.580 75.320 ;
        RECT 76.110 75.000 76.370 75.320 ;
        RECT 76.700 75.000 76.960 75.320 ;
        RECT 77.505 75.245 77.735 76.555 ;
        RECT 78.345 75.245 78.515 77.185 ;
        RECT 77.505 75.075 78.515 75.245 ;
        RECT 78.660 75.075 79.015 77.185 ;
        RECT 79.385 77.185 81.395 77.365 ;
        RECT 82.330 77.460 82.570 77.690 ;
        RECT 86.485 77.685 87.895 77.925 ;
        RECT 82.330 77.360 84.235 77.460 ;
        RECT 86.485 77.425 86.725 77.685 ;
        RECT 84.820 77.365 86.725 77.425 ;
        RECT 82.330 77.220 84.340 77.360 ;
        RECT 83.670 77.185 84.340 77.220 ;
        RECT 79.385 75.080 79.740 77.185 ;
        RECT 80.660 75.320 80.890 76.555 ;
        RECT 81.450 75.320 81.680 76.555 ;
        RECT 82.040 75.320 82.270 76.555 ;
        RECT 75.335 74.110 75.565 75.000 ;
        RECT 76.125 74.110 76.355 75.000 ;
        RECT 76.715 74.110 76.945 75.000 ;
        RECT 77.505 74.110 77.735 75.075 ;
        RECT 80.645 75.000 80.905 75.320 ;
        RECT 81.435 75.000 81.695 75.320 ;
        RECT 82.025 75.000 82.285 75.320 ;
        RECT 82.830 75.245 83.060 76.555 ;
        RECT 83.670 75.245 83.840 77.185 ;
        RECT 82.830 75.075 83.840 75.245 ;
        RECT 83.985 75.075 84.340 77.185 ;
        RECT 84.720 77.185 86.725 77.365 ;
        RECT 87.655 77.460 87.895 77.685 ;
        RECT 91.815 77.690 93.230 77.930 ;
        RECT 87.655 77.360 89.570 77.460 ;
        RECT 91.815 77.425 92.055 77.690 ;
        RECT 90.145 77.365 92.055 77.425 ;
        RECT 87.655 77.220 89.675 77.360 ;
        RECT 89.005 77.185 89.675 77.220 ;
        RECT 84.720 75.080 85.075 77.185 ;
        RECT 85.995 75.320 86.225 76.555 ;
        RECT 86.785 75.320 87.015 76.555 ;
        RECT 87.375 75.320 87.605 76.555 ;
        RECT 80.660 74.110 80.890 75.000 ;
        RECT 81.450 74.110 81.680 75.000 ;
        RECT 82.040 74.110 82.270 75.000 ;
        RECT 82.830 74.110 83.060 75.075 ;
        RECT 85.980 75.000 86.240 75.320 ;
        RECT 86.770 75.000 87.030 75.320 ;
        RECT 87.360 75.000 87.620 75.320 ;
        RECT 88.165 75.245 88.395 76.555 ;
        RECT 89.005 75.245 89.175 77.185 ;
        RECT 88.165 75.075 89.175 75.245 ;
        RECT 89.320 75.075 89.675 77.185 ;
        RECT 90.045 77.185 92.055 77.365 ;
        RECT 92.990 77.460 93.230 77.690 ;
        RECT 97.145 77.685 98.555 77.925 ;
        RECT 92.990 77.360 94.895 77.460 ;
        RECT 97.145 77.425 97.385 77.685 ;
        RECT 95.480 77.365 97.385 77.425 ;
        RECT 92.990 77.220 95.000 77.360 ;
        RECT 94.330 77.185 95.000 77.220 ;
        RECT 90.045 75.080 90.400 77.185 ;
        RECT 91.320 75.320 91.550 76.555 ;
        RECT 92.110 75.320 92.340 76.555 ;
        RECT 92.700 75.320 92.930 76.555 ;
        RECT 85.995 74.110 86.225 75.000 ;
        RECT 86.785 74.110 87.015 75.000 ;
        RECT 87.375 74.110 87.605 75.000 ;
        RECT 88.165 74.110 88.395 75.075 ;
        RECT 91.305 75.000 91.565 75.320 ;
        RECT 92.095 75.000 92.355 75.320 ;
        RECT 92.685 75.000 92.945 75.320 ;
        RECT 93.490 75.245 93.720 76.555 ;
        RECT 94.330 75.245 94.500 77.185 ;
        RECT 93.490 75.075 94.500 75.245 ;
        RECT 94.645 75.075 95.000 77.185 ;
        RECT 95.380 77.185 97.385 77.365 ;
        RECT 98.315 77.460 98.555 77.685 ;
        RECT 102.475 77.690 103.890 77.930 ;
        RECT 98.315 77.360 100.230 77.460 ;
        RECT 102.475 77.425 102.715 77.690 ;
        RECT 100.805 77.365 102.715 77.425 ;
        RECT 98.315 77.220 100.335 77.360 ;
        RECT 99.665 77.185 100.335 77.220 ;
        RECT 95.380 75.080 95.735 77.185 ;
        RECT 96.655 75.320 96.885 76.555 ;
        RECT 97.445 75.320 97.675 76.555 ;
        RECT 98.035 75.320 98.265 76.555 ;
        RECT 91.320 74.110 91.550 75.000 ;
        RECT 92.110 74.110 92.340 75.000 ;
        RECT 92.700 74.110 92.930 75.000 ;
        RECT 93.490 74.110 93.720 75.075 ;
        RECT 96.640 75.000 96.900 75.320 ;
        RECT 97.430 75.000 97.690 75.320 ;
        RECT 98.020 75.000 98.280 75.320 ;
        RECT 98.825 75.245 99.055 76.555 ;
        RECT 99.665 75.245 99.835 77.185 ;
        RECT 98.825 75.075 99.835 75.245 ;
        RECT 99.980 75.075 100.335 77.185 ;
        RECT 100.705 77.185 102.715 77.365 ;
        RECT 103.650 77.460 103.890 77.690 ;
        RECT 107.805 77.685 109.215 77.925 ;
        RECT 103.650 77.360 105.555 77.460 ;
        RECT 107.805 77.425 108.045 77.685 ;
        RECT 106.140 77.365 108.045 77.425 ;
        RECT 103.650 77.220 105.660 77.360 ;
        RECT 104.990 77.185 105.660 77.220 ;
        RECT 100.705 75.080 101.060 77.185 ;
        RECT 101.980 75.320 102.210 76.555 ;
        RECT 102.770 75.320 103.000 76.555 ;
        RECT 103.360 75.320 103.590 76.555 ;
        RECT 96.655 74.110 96.885 75.000 ;
        RECT 97.445 74.110 97.675 75.000 ;
        RECT 98.035 74.110 98.265 75.000 ;
        RECT 98.825 74.110 99.055 75.075 ;
        RECT 101.965 75.000 102.225 75.320 ;
        RECT 102.755 75.000 103.015 75.320 ;
        RECT 103.345 75.000 103.605 75.320 ;
        RECT 104.150 75.245 104.380 76.555 ;
        RECT 104.990 75.245 105.160 77.185 ;
        RECT 104.150 75.075 105.160 75.245 ;
        RECT 105.305 75.075 105.660 77.185 ;
        RECT 106.040 77.185 108.045 77.365 ;
        RECT 108.975 77.460 109.215 77.685 ;
        RECT 113.135 77.690 114.550 77.930 ;
        RECT 108.975 77.360 110.890 77.460 ;
        RECT 113.135 77.425 113.375 77.690 ;
        RECT 111.465 77.365 113.375 77.425 ;
        RECT 108.975 77.220 110.995 77.360 ;
        RECT 110.325 77.185 110.995 77.220 ;
        RECT 106.040 75.080 106.395 77.185 ;
        RECT 107.315 75.320 107.545 76.555 ;
        RECT 108.105 75.320 108.335 76.555 ;
        RECT 108.695 75.320 108.925 76.555 ;
        RECT 101.980 74.110 102.210 75.000 ;
        RECT 102.770 74.110 103.000 75.000 ;
        RECT 103.360 74.110 103.590 75.000 ;
        RECT 104.150 74.110 104.380 75.075 ;
        RECT 107.300 75.000 107.560 75.320 ;
        RECT 108.090 75.000 108.350 75.320 ;
        RECT 108.680 75.000 108.940 75.320 ;
        RECT 109.485 75.245 109.715 76.555 ;
        RECT 110.325 75.245 110.495 77.185 ;
        RECT 109.485 75.075 110.495 75.245 ;
        RECT 110.640 75.075 110.995 77.185 ;
        RECT 111.365 77.185 113.375 77.365 ;
        RECT 114.310 77.460 114.550 77.690 ;
        RECT 118.465 77.685 119.875 77.925 ;
        RECT 114.310 77.360 116.215 77.460 ;
        RECT 118.465 77.425 118.705 77.685 ;
        RECT 116.800 77.365 118.705 77.425 ;
        RECT 114.310 77.220 116.320 77.360 ;
        RECT 115.650 77.185 116.320 77.220 ;
        RECT 111.365 75.080 111.720 77.185 ;
        RECT 112.640 75.320 112.870 76.555 ;
        RECT 113.430 75.320 113.660 76.555 ;
        RECT 114.020 75.320 114.250 76.555 ;
        RECT 107.315 74.110 107.545 75.000 ;
        RECT 108.105 74.110 108.335 75.000 ;
        RECT 108.695 74.110 108.925 75.000 ;
        RECT 109.485 74.110 109.715 75.075 ;
        RECT 112.625 75.000 112.885 75.320 ;
        RECT 113.415 75.000 113.675 75.320 ;
        RECT 114.005 75.000 114.265 75.320 ;
        RECT 114.810 75.245 115.040 76.555 ;
        RECT 115.650 75.245 115.820 77.185 ;
        RECT 114.810 75.075 115.820 75.245 ;
        RECT 115.965 75.075 116.320 77.185 ;
        RECT 116.700 77.185 118.705 77.365 ;
        RECT 119.635 77.460 119.875 77.685 ;
        RECT 123.240 77.705 125.790 77.970 ;
        RECT 123.240 77.500 123.575 77.705 ;
        RECT 119.635 77.360 121.550 77.460 ;
        RECT 122.075 77.380 123.575 77.500 ;
        RECT 119.635 77.220 121.655 77.360 ;
        RECT 120.985 77.185 121.655 77.220 ;
        RECT 116.700 75.080 117.055 77.185 ;
        RECT 117.975 75.320 118.205 76.555 ;
        RECT 118.765 75.320 118.995 76.555 ;
        RECT 119.355 75.320 119.585 76.555 ;
        RECT 112.640 74.110 112.870 75.000 ;
        RECT 113.430 74.110 113.660 75.000 ;
        RECT 114.020 74.110 114.250 75.000 ;
        RECT 114.810 74.110 115.040 75.075 ;
        RECT 117.960 75.000 118.220 75.320 ;
        RECT 118.750 75.000 119.010 75.320 ;
        RECT 119.340 75.000 119.600 75.320 ;
        RECT 120.145 75.245 120.375 76.555 ;
        RECT 120.985 75.245 121.155 77.185 ;
        RECT 120.145 75.075 121.155 75.245 ;
        RECT 121.300 75.075 121.655 77.185 ;
        RECT 122.025 77.185 123.575 77.380 ;
        RECT 125.455 77.460 125.790 77.705 ;
        RECT 125.455 77.380 126.875 77.460 ;
        RECT 125.455 77.185 126.980 77.380 ;
        RECT 122.025 77.165 122.425 77.185 ;
        RECT 122.025 75.095 122.380 77.165 ;
        RECT 123.300 75.320 123.530 76.555 ;
        RECT 124.090 75.320 124.320 76.555 ;
        RECT 124.680 75.320 124.910 76.555 ;
        RECT 117.975 74.110 118.205 75.000 ;
        RECT 118.765 74.110 118.995 75.000 ;
        RECT 119.355 74.110 119.585 75.000 ;
        RECT 120.145 74.110 120.375 75.075 ;
        RECT 123.285 75.000 123.545 75.320 ;
        RECT 124.075 75.000 124.335 75.320 ;
        RECT 124.665 75.000 124.925 75.320 ;
        RECT 125.470 75.245 125.700 76.555 ;
        RECT 126.310 75.245 126.480 77.185 ;
        RECT 125.470 75.075 126.480 75.245 ;
        RECT 126.625 75.095 126.980 77.185 ;
        RECT 123.300 74.110 123.530 75.000 ;
        RECT 124.090 74.110 124.320 75.000 ;
        RECT 124.680 74.110 124.910 75.000 ;
        RECT 125.470 74.110 125.700 75.075 ;
        RECT 31.420 69.925 31.775 72.135 ;
        RECT 32.695 72.055 32.925 73.020 ;
        RECT 33.485 72.145 33.715 73.020 ;
        RECT 34.075 72.145 34.305 73.020 ;
        RECT 34.865 72.145 35.095 73.020 ;
        RECT 31.915 71.885 32.925 72.055 ;
        RECT 31.915 69.925 32.085 71.885 ;
        RECT 32.695 70.575 32.925 71.885 ;
        RECT 33.470 71.825 33.730 72.145 ;
        RECT 34.060 71.825 34.320 72.145 ;
        RECT 34.850 71.825 35.110 72.145 ;
        RECT 33.485 70.575 33.715 71.825 ;
        RECT 34.075 70.575 34.305 71.825 ;
        RECT 34.865 70.575 35.095 71.825 ;
        RECT 36.020 69.925 36.375 72.135 ;
        RECT 31.420 69.650 32.085 69.925 ;
        RECT 35.705 69.650 36.375 69.925 ;
        RECT 31.420 67.560 31.775 69.650 ;
        RECT 32.695 67.785 32.925 69.020 ;
        RECT 33.485 67.785 33.715 69.020 ;
        RECT 34.075 67.785 34.305 69.020 ;
        RECT 31.510 67.540 31.770 67.560 ;
        RECT 32.680 67.465 32.940 67.785 ;
        RECT 33.470 67.465 33.730 67.785 ;
        RECT 34.060 67.465 34.320 67.785 ;
        RECT 34.865 67.710 35.095 69.020 ;
        RECT 35.705 67.710 35.875 69.650 ;
        RECT 36.020 67.855 36.375 69.650 ;
        RECT 34.865 67.540 35.875 67.710 ;
        RECT 36.015 67.560 36.375 67.855 ;
        RECT 36.745 69.925 37.100 72.120 ;
        RECT 38.020 72.055 38.250 73.020 ;
        RECT 38.810 72.145 39.040 73.020 ;
        RECT 39.400 72.145 39.630 73.020 ;
        RECT 40.190 72.145 40.420 73.020 ;
        RECT 37.240 71.885 38.250 72.055 ;
        RECT 37.240 69.925 37.410 71.885 ;
        RECT 38.020 70.575 38.250 71.885 ;
        RECT 38.795 71.825 39.055 72.145 ;
        RECT 39.385 71.825 39.645 72.145 ;
        RECT 40.175 71.825 40.435 72.145 ;
        RECT 38.810 70.575 39.040 71.825 ;
        RECT 39.400 70.575 39.630 71.825 ;
        RECT 40.190 70.575 40.420 71.825 ;
        RECT 41.345 69.925 41.700 72.115 ;
        RECT 36.745 69.650 37.410 69.925 ;
        RECT 41.030 69.650 41.700 69.925 ;
        RECT 32.695 66.575 32.925 67.465 ;
        RECT 33.485 66.575 33.715 67.465 ;
        RECT 34.075 66.575 34.305 67.465 ;
        RECT 34.865 66.575 35.095 67.540 ;
        RECT 36.015 67.535 36.275 67.560 ;
        RECT 36.745 67.545 37.100 69.650 ;
        RECT 37.520 69.225 38.760 69.455 ;
        RECT 39.680 69.225 40.870 69.455 ;
        RECT 37.520 68.800 37.780 69.225 ;
        RECT 38.020 67.785 38.250 69.020 ;
        RECT 38.810 67.785 39.040 69.020 ;
        RECT 39.400 67.785 39.630 69.020 ;
        RECT 38.005 67.465 38.265 67.785 ;
        RECT 38.795 67.465 39.055 67.785 ;
        RECT 39.385 67.465 39.645 67.785 ;
        RECT 40.190 67.710 40.420 69.020 ;
        RECT 40.610 67.850 40.870 69.225 ;
        RECT 41.030 67.710 41.200 69.650 ;
        RECT 41.345 69.140 41.700 69.650 ;
        RECT 41.340 68.350 41.700 69.140 ;
        RECT 40.190 67.540 41.200 67.710 ;
        RECT 41.345 67.540 41.700 68.350 ;
        RECT 42.080 69.925 42.435 72.120 ;
        RECT 43.355 72.055 43.585 73.020 ;
        RECT 44.145 72.145 44.375 73.020 ;
        RECT 44.735 72.145 44.965 73.020 ;
        RECT 45.525 72.145 45.755 73.020 ;
        RECT 42.575 71.885 43.585 72.055 ;
        RECT 42.575 69.925 42.745 71.885 ;
        RECT 43.355 70.575 43.585 71.885 ;
        RECT 44.130 71.825 44.390 72.145 ;
        RECT 44.720 71.825 44.980 72.145 ;
        RECT 45.510 71.825 45.770 72.145 ;
        RECT 44.145 70.575 44.375 71.825 ;
        RECT 44.735 70.575 44.965 71.825 ;
        RECT 45.525 70.575 45.755 71.825 ;
        RECT 46.680 69.925 47.035 72.115 ;
        RECT 42.080 69.650 42.745 69.925 ;
        RECT 46.365 69.650 47.035 69.925 ;
        RECT 42.080 67.545 42.435 69.650 ;
        RECT 42.855 69.225 44.095 69.455 ;
        RECT 45.015 69.225 46.205 69.455 ;
        RECT 42.855 68.800 43.115 69.225 ;
        RECT 43.355 67.785 43.585 69.020 ;
        RECT 44.145 67.785 44.375 69.020 ;
        RECT 44.735 67.785 44.965 69.020 ;
        RECT 37.520 66.415 37.780 67.295 ;
        RECT 38.020 66.575 38.250 67.465 ;
        RECT 38.810 66.575 39.040 67.465 ;
        RECT 39.400 66.575 39.630 67.465 ;
        RECT 40.190 66.575 40.420 67.540 ;
        RECT 43.340 67.465 43.600 67.785 ;
        RECT 44.130 67.465 44.390 67.785 ;
        RECT 44.720 67.465 44.980 67.785 ;
        RECT 45.525 67.710 45.755 69.020 ;
        RECT 45.945 67.850 46.205 69.225 ;
        RECT 46.365 67.710 46.535 69.650 ;
        RECT 46.680 69.140 47.035 69.650 ;
        RECT 46.675 68.350 47.035 69.140 ;
        RECT 45.525 67.540 46.535 67.710 ;
        RECT 46.680 67.540 47.035 68.350 ;
        RECT 47.405 69.925 47.760 72.120 ;
        RECT 48.680 72.055 48.910 73.020 ;
        RECT 49.470 72.145 49.700 73.020 ;
        RECT 50.060 72.145 50.290 73.020 ;
        RECT 50.850 72.145 51.080 73.020 ;
        RECT 47.900 71.885 48.910 72.055 ;
        RECT 47.900 69.925 48.070 71.885 ;
        RECT 48.680 70.575 48.910 71.885 ;
        RECT 49.455 71.825 49.715 72.145 ;
        RECT 50.045 71.825 50.305 72.145 ;
        RECT 50.835 71.825 51.095 72.145 ;
        RECT 49.470 70.575 49.700 71.825 ;
        RECT 50.060 70.575 50.290 71.825 ;
        RECT 50.850 70.575 51.080 71.825 ;
        RECT 52.005 69.925 52.360 72.115 ;
        RECT 47.405 69.650 48.070 69.925 ;
        RECT 51.690 69.650 52.360 69.925 ;
        RECT 47.405 67.545 47.760 69.650 ;
        RECT 48.180 69.225 49.420 69.455 ;
        RECT 50.340 69.225 51.530 69.455 ;
        RECT 48.180 68.800 48.440 69.225 ;
        RECT 48.680 67.785 48.910 69.020 ;
        RECT 49.470 67.785 49.700 69.020 ;
        RECT 50.060 67.785 50.290 69.020 ;
        RECT 40.660 66.415 40.920 67.205 ;
        RECT 37.520 66.185 38.760 66.415 ;
        RECT 39.680 66.185 40.920 66.415 ;
        RECT 42.855 66.415 43.115 67.295 ;
        RECT 43.355 66.575 43.585 67.465 ;
        RECT 44.145 66.575 44.375 67.465 ;
        RECT 44.735 66.575 44.965 67.465 ;
        RECT 45.525 66.575 45.755 67.540 ;
        RECT 48.665 67.465 48.925 67.785 ;
        RECT 49.455 67.465 49.715 67.785 ;
        RECT 50.045 67.465 50.305 67.785 ;
        RECT 50.850 67.710 51.080 69.020 ;
        RECT 51.270 67.850 51.530 69.225 ;
        RECT 51.690 67.710 51.860 69.650 ;
        RECT 52.005 69.140 52.360 69.650 ;
        RECT 52.000 68.350 52.360 69.140 ;
        RECT 50.850 67.540 51.860 67.710 ;
        RECT 52.005 67.540 52.360 68.350 ;
        RECT 52.740 69.925 53.095 72.120 ;
        RECT 54.015 72.055 54.245 73.020 ;
        RECT 54.805 72.145 55.035 73.020 ;
        RECT 55.395 72.145 55.625 73.020 ;
        RECT 56.185 72.145 56.415 73.020 ;
        RECT 53.235 71.885 54.245 72.055 ;
        RECT 53.235 69.925 53.405 71.885 ;
        RECT 54.015 70.575 54.245 71.885 ;
        RECT 54.790 71.825 55.050 72.145 ;
        RECT 55.380 71.825 55.640 72.145 ;
        RECT 56.170 71.825 56.430 72.145 ;
        RECT 54.805 70.575 55.035 71.825 ;
        RECT 55.395 70.575 55.625 71.825 ;
        RECT 56.185 70.575 56.415 71.825 ;
        RECT 57.340 69.925 57.695 72.115 ;
        RECT 52.740 69.650 53.405 69.925 ;
        RECT 57.025 69.650 57.695 69.925 ;
        RECT 52.740 67.545 53.095 69.650 ;
        RECT 53.515 69.225 54.755 69.455 ;
        RECT 55.675 69.225 56.865 69.455 ;
        RECT 53.515 68.800 53.775 69.225 ;
        RECT 54.805 67.785 55.035 69.020 ;
        RECT 55.395 67.785 55.625 69.020 ;
        RECT 45.995 66.415 46.255 67.205 ;
        RECT 42.855 66.185 44.095 66.415 ;
        RECT 45.015 66.185 46.255 66.415 ;
        RECT 48.180 66.415 48.440 67.295 ;
        RECT 48.680 66.575 48.910 67.465 ;
        RECT 49.470 66.575 49.700 67.465 ;
        RECT 50.060 66.575 50.290 67.465 ;
        RECT 50.850 66.575 51.080 67.540 ;
        RECT 54.790 67.465 55.050 67.785 ;
        RECT 55.380 67.465 55.640 67.785 ;
        RECT 56.185 67.710 56.415 69.020 ;
        RECT 56.605 67.850 56.865 69.225 ;
        RECT 57.025 67.710 57.195 69.650 ;
        RECT 57.340 69.140 57.695 69.650 ;
        RECT 57.335 68.350 57.695 69.140 ;
        RECT 56.185 67.540 57.195 67.710 ;
        RECT 57.340 67.540 57.695 68.350 ;
        RECT 58.065 69.925 58.420 72.120 ;
        RECT 59.340 72.055 59.570 73.020 ;
        RECT 60.130 72.145 60.360 73.020 ;
        RECT 60.720 72.145 60.950 73.020 ;
        RECT 61.510 72.145 61.740 73.020 ;
        RECT 58.560 71.885 59.570 72.055 ;
        RECT 58.560 69.925 58.730 71.885 ;
        RECT 59.340 70.575 59.570 71.885 ;
        RECT 60.115 71.825 60.375 72.145 ;
        RECT 60.705 71.825 60.965 72.145 ;
        RECT 61.495 71.825 61.755 72.145 ;
        RECT 60.130 70.575 60.360 71.825 ;
        RECT 60.720 70.575 60.950 71.825 ;
        RECT 61.510 70.575 61.740 71.825 ;
        RECT 62.665 69.925 63.020 72.115 ;
        RECT 58.065 69.650 58.730 69.925 ;
        RECT 62.350 69.650 63.020 69.925 ;
        RECT 58.065 67.545 58.420 69.650 ;
        RECT 58.840 69.225 60.080 69.455 ;
        RECT 61.000 69.225 62.190 69.455 ;
        RECT 58.840 68.800 59.100 69.225 ;
        RECT 59.340 67.785 59.570 69.020 ;
        RECT 60.130 67.785 60.360 69.020 ;
        RECT 60.720 67.785 60.950 69.020 ;
        RECT 51.320 66.415 51.580 67.205 ;
        RECT 48.180 66.185 49.420 66.415 ;
        RECT 50.340 66.185 51.580 66.415 ;
        RECT 53.515 66.415 53.775 67.295 ;
        RECT 54.805 66.575 55.035 67.465 ;
        RECT 55.395 66.575 55.625 67.465 ;
        RECT 56.185 66.575 56.415 67.540 ;
        RECT 59.325 67.465 59.585 67.785 ;
        RECT 60.115 67.465 60.375 67.785 ;
        RECT 60.705 67.465 60.965 67.785 ;
        RECT 61.510 67.710 61.740 69.020 ;
        RECT 61.930 67.850 62.190 69.225 ;
        RECT 62.350 67.710 62.520 69.650 ;
        RECT 62.665 69.140 63.020 69.650 ;
        RECT 62.660 68.350 63.020 69.140 ;
        RECT 61.510 67.540 62.520 67.710 ;
        RECT 62.665 67.540 63.020 68.350 ;
        RECT 63.400 69.925 63.755 72.120 ;
        RECT 64.675 72.055 64.905 73.020 ;
        RECT 65.465 72.145 65.695 73.020 ;
        RECT 66.055 72.145 66.285 73.020 ;
        RECT 66.845 72.145 67.075 73.020 ;
        RECT 63.895 71.885 64.905 72.055 ;
        RECT 63.895 69.925 64.065 71.885 ;
        RECT 64.675 70.575 64.905 71.885 ;
        RECT 65.450 71.825 65.710 72.145 ;
        RECT 66.040 71.825 66.300 72.145 ;
        RECT 66.830 71.825 67.090 72.145 ;
        RECT 65.465 70.575 65.695 71.825 ;
        RECT 66.055 70.575 66.285 71.825 ;
        RECT 66.845 70.575 67.075 71.825 ;
        RECT 68.000 69.925 68.355 72.115 ;
        RECT 63.400 69.650 64.065 69.925 ;
        RECT 67.685 69.650 68.355 69.925 ;
        RECT 63.400 67.545 63.755 69.650 ;
        RECT 64.175 69.225 65.415 69.455 ;
        RECT 66.335 69.225 67.525 69.455 ;
        RECT 64.175 68.800 64.435 69.225 ;
        RECT 64.675 67.785 64.905 69.020 ;
        RECT 65.465 67.785 65.695 69.020 ;
        RECT 66.055 67.785 66.285 69.020 ;
        RECT 56.655 66.415 56.915 67.205 ;
        RECT 53.515 66.185 54.755 66.415 ;
        RECT 55.675 66.185 56.915 66.415 ;
        RECT 58.840 66.415 59.100 67.295 ;
        RECT 59.340 66.575 59.570 67.465 ;
        RECT 60.130 66.575 60.360 67.465 ;
        RECT 60.720 66.575 60.950 67.465 ;
        RECT 61.510 66.575 61.740 67.540 ;
        RECT 64.660 67.465 64.920 67.785 ;
        RECT 65.450 67.465 65.710 67.785 ;
        RECT 66.040 67.465 66.300 67.785 ;
        RECT 66.845 67.710 67.075 69.020 ;
        RECT 67.265 67.850 67.525 69.225 ;
        RECT 67.685 67.710 67.855 69.650 ;
        RECT 68.000 69.140 68.355 69.650 ;
        RECT 67.995 68.350 68.355 69.140 ;
        RECT 66.845 67.540 67.855 67.710 ;
        RECT 68.000 67.540 68.355 68.350 ;
        RECT 68.725 69.925 69.080 72.120 ;
        RECT 70.000 72.055 70.230 73.020 ;
        RECT 70.790 72.145 71.020 73.020 ;
        RECT 71.380 72.145 71.610 73.020 ;
        RECT 72.170 72.145 72.400 73.020 ;
        RECT 69.220 71.885 70.230 72.055 ;
        RECT 69.220 69.925 69.390 71.885 ;
        RECT 70.000 70.575 70.230 71.885 ;
        RECT 70.775 71.825 71.035 72.145 ;
        RECT 71.365 71.825 71.625 72.145 ;
        RECT 72.155 71.825 72.415 72.145 ;
        RECT 70.790 70.575 71.020 71.825 ;
        RECT 71.380 70.575 71.610 71.825 ;
        RECT 72.170 70.575 72.400 71.825 ;
        RECT 73.325 69.925 73.680 72.115 ;
        RECT 68.725 69.650 69.390 69.925 ;
        RECT 73.010 69.650 73.680 69.925 ;
        RECT 68.725 67.545 69.080 69.650 ;
        RECT 69.500 69.225 70.740 69.455 ;
        RECT 71.660 69.225 72.850 69.455 ;
        RECT 69.500 68.800 69.760 69.225 ;
        RECT 70.000 67.785 70.230 69.020 ;
        RECT 70.790 67.785 71.020 69.020 ;
        RECT 71.380 67.785 71.610 69.020 ;
        RECT 61.980 66.415 62.240 67.205 ;
        RECT 58.840 66.185 60.080 66.415 ;
        RECT 61.000 66.185 62.240 66.415 ;
        RECT 64.175 66.415 64.435 67.295 ;
        RECT 64.675 66.575 64.905 67.465 ;
        RECT 65.465 66.575 65.695 67.465 ;
        RECT 66.055 66.575 66.285 67.465 ;
        RECT 66.845 66.575 67.075 67.540 ;
        RECT 69.985 67.465 70.245 67.785 ;
        RECT 70.775 67.465 71.035 67.785 ;
        RECT 71.365 67.465 71.625 67.785 ;
        RECT 72.170 67.710 72.400 69.020 ;
        RECT 72.590 67.850 72.850 69.225 ;
        RECT 73.010 67.710 73.180 69.650 ;
        RECT 73.325 69.140 73.680 69.650 ;
        RECT 73.320 68.350 73.680 69.140 ;
        RECT 72.170 67.540 73.180 67.710 ;
        RECT 73.325 67.540 73.680 68.350 ;
        RECT 74.060 69.925 74.415 72.120 ;
        RECT 75.335 72.055 75.565 73.020 ;
        RECT 76.125 72.145 76.355 73.020 ;
        RECT 76.715 72.145 76.945 73.020 ;
        RECT 77.505 72.145 77.735 73.020 ;
        RECT 74.555 71.885 75.565 72.055 ;
        RECT 74.555 69.925 74.725 71.885 ;
        RECT 75.335 70.575 75.565 71.885 ;
        RECT 76.110 71.825 76.370 72.145 ;
        RECT 76.700 71.825 76.960 72.145 ;
        RECT 77.490 71.825 77.750 72.145 ;
        RECT 76.125 70.575 76.355 71.825 ;
        RECT 76.715 70.575 76.945 71.825 ;
        RECT 77.505 70.575 77.735 71.825 ;
        RECT 78.660 69.925 79.015 72.115 ;
        RECT 74.060 69.650 74.725 69.925 ;
        RECT 78.345 69.650 79.015 69.925 ;
        RECT 74.060 67.545 74.415 69.650 ;
        RECT 76.995 69.225 78.185 69.455 ;
        RECT 75.335 67.785 75.565 69.020 ;
        RECT 76.125 67.785 76.355 69.020 ;
        RECT 76.715 67.785 76.945 69.020 ;
        RECT 67.315 66.415 67.575 67.205 ;
        RECT 64.175 66.185 65.415 66.415 ;
        RECT 66.335 66.185 67.575 66.415 ;
        RECT 69.500 66.415 69.760 67.295 ;
        RECT 70.000 66.575 70.230 67.465 ;
        RECT 70.790 66.575 71.020 67.465 ;
        RECT 71.380 66.575 71.610 67.465 ;
        RECT 72.170 66.575 72.400 67.540 ;
        RECT 75.320 67.465 75.580 67.785 ;
        RECT 76.110 67.465 76.370 67.785 ;
        RECT 76.700 67.465 76.960 67.785 ;
        RECT 77.505 67.710 77.735 69.020 ;
        RECT 77.925 67.850 78.185 69.225 ;
        RECT 78.345 67.710 78.515 69.650 ;
        RECT 78.660 69.140 79.015 69.650 ;
        RECT 78.655 68.350 79.015 69.140 ;
        RECT 77.505 67.540 78.515 67.710 ;
        RECT 78.660 67.540 79.015 68.350 ;
        RECT 79.385 69.925 79.740 72.120 ;
        RECT 80.660 72.055 80.890 73.020 ;
        RECT 81.450 72.145 81.680 73.020 ;
        RECT 82.040 72.145 82.270 73.020 ;
        RECT 82.830 72.145 83.060 73.020 ;
        RECT 79.880 71.885 80.890 72.055 ;
        RECT 79.880 69.925 80.050 71.885 ;
        RECT 80.660 70.575 80.890 71.885 ;
        RECT 81.435 71.825 81.695 72.145 ;
        RECT 82.025 71.825 82.285 72.145 ;
        RECT 82.815 71.825 83.075 72.145 ;
        RECT 81.450 70.575 81.680 71.825 ;
        RECT 82.040 70.575 82.270 71.825 ;
        RECT 82.830 70.575 83.060 71.825 ;
        RECT 83.985 69.925 84.340 72.115 ;
        RECT 79.385 69.650 80.050 69.925 ;
        RECT 83.670 69.650 84.340 69.925 ;
        RECT 79.385 67.545 79.740 69.650 ;
        RECT 80.160 69.225 81.400 69.455 ;
        RECT 82.320 69.225 83.510 69.455 ;
        RECT 80.160 68.800 80.420 69.225 ;
        RECT 80.660 67.785 80.890 69.020 ;
        RECT 81.450 67.785 81.680 69.020 ;
        RECT 82.040 67.785 82.270 69.020 ;
        RECT 72.640 66.415 72.900 67.205 ;
        RECT 75.335 66.575 75.565 67.465 ;
        RECT 76.125 66.575 76.355 67.465 ;
        RECT 76.715 66.575 76.945 67.465 ;
        RECT 77.505 66.575 77.735 67.540 ;
        RECT 80.645 67.465 80.905 67.785 ;
        RECT 81.435 67.465 81.695 67.785 ;
        RECT 82.025 67.465 82.285 67.785 ;
        RECT 82.830 67.710 83.060 69.020 ;
        RECT 83.250 67.850 83.510 69.225 ;
        RECT 83.670 67.710 83.840 69.650 ;
        RECT 83.985 69.140 84.340 69.650 ;
        RECT 83.980 68.350 84.340 69.140 ;
        RECT 82.830 67.540 83.840 67.710 ;
        RECT 83.985 67.540 84.340 68.350 ;
        RECT 84.720 69.925 85.075 72.120 ;
        RECT 85.995 72.055 86.225 73.020 ;
        RECT 86.785 72.145 87.015 73.020 ;
        RECT 87.375 72.145 87.605 73.020 ;
        RECT 88.165 72.145 88.395 73.020 ;
        RECT 85.215 71.885 86.225 72.055 ;
        RECT 85.215 69.925 85.385 71.885 ;
        RECT 85.995 70.575 86.225 71.885 ;
        RECT 86.770 71.825 87.030 72.145 ;
        RECT 87.360 71.825 87.620 72.145 ;
        RECT 88.150 71.825 88.410 72.145 ;
        RECT 86.785 70.575 87.015 71.825 ;
        RECT 87.375 70.575 87.605 71.825 ;
        RECT 88.165 70.575 88.395 71.825 ;
        RECT 89.320 69.925 89.675 72.115 ;
        RECT 84.720 69.650 85.385 69.925 ;
        RECT 89.005 69.650 89.675 69.925 ;
        RECT 84.720 67.545 85.075 69.650 ;
        RECT 85.495 69.225 86.735 69.455 ;
        RECT 87.655 69.225 88.845 69.455 ;
        RECT 85.495 68.800 85.755 69.225 ;
        RECT 85.995 67.785 86.225 69.020 ;
        RECT 86.785 67.785 87.015 69.020 ;
        RECT 87.375 67.785 87.605 69.020 ;
        RECT 77.975 66.415 78.235 67.205 ;
        RECT 69.500 66.185 70.740 66.415 ;
        RECT 71.660 66.185 72.900 66.415 ;
        RECT 76.995 66.185 78.235 66.415 ;
        RECT 80.160 66.415 80.420 67.295 ;
        RECT 80.660 66.575 80.890 67.465 ;
        RECT 81.450 66.575 81.680 67.465 ;
        RECT 82.040 66.575 82.270 67.465 ;
        RECT 82.830 66.575 83.060 67.540 ;
        RECT 85.980 67.465 86.240 67.785 ;
        RECT 86.770 67.465 87.030 67.785 ;
        RECT 87.360 67.465 87.620 67.785 ;
        RECT 88.165 67.710 88.395 69.020 ;
        RECT 88.585 67.850 88.845 69.225 ;
        RECT 89.005 67.710 89.175 69.650 ;
        RECT 89.320 69.140 89.675 69.650 ;
        RECT 89.315 68.350 89.675 69.140 ;
        RECT 88.165 67.540 89.175 67.710 ;
        RECT 89.320 67.540 89.675 68.350 ;
        RECT 90.045 69.925 90.400 72.120 ;
        RECT 91.320 72.055 91.550 73.020 ;
        RECT 92.110 72.145 92.340 73.020 ;
        RECT 92.700 72.145 92.930 73.020 ;
        RECT 93.490 72.145 93.720 73.020 ;
        RECT 90.540 71.885 91.550 72.055 ;
        RECT 90.540 69.925 90.710 71.885 ;
        RECT 91.320 70.575 91.550 71.885 ;
        RECT 92.095 71.825 92.355 72.145 ;
        RECT 92.685 71.825 92.945 72.145 ;
        RECT 93.475 71.825 93.735 72.145 ;
        RECT 92.110 70.575 92.340 71.825 ;
        RECT 92.700 70.575 92.930 71.825 ;
        RECT 93.490 70.575 93.720 71.825 ;
        RECT 94.645 69.925 95.000 72.115 ;
        RECT 90.045 69.650 90.710 69.925 ;
        RECT 94.330 69.650 95.000 69.925 ;
        RECT 90.045 67.545 90.400 69.650 ;
        RECT 90.820 69.225 92.060 69.455 ;
        RECT 92.980 69.225 94.170 69.455 ;
        RECT 90.820 68.800 91.080 69.225 ;
        RECT 91.320 67.785 91.550 69.020 ;
        RECT 92.110 67.785 92.340 69.020 ;
        RECT 92.700 67.785 92.930 69.020 ;
        RECT 83.300 66.415 83.560 67.205 ;
        RECT 80.160 66.185 81.400 66.415 ;
        RECT 82.320 66.185 83.560 66.415 ;
        RECT 85.495 66.415 85.755 67.295 ;
        RECT 85.995 66.575 86.225 67.465 ;
        RECT 86.785 66.575 87.015 67.465 ;
        RECT 87.375 66.575 87.605 67.465 ;
        RECT 88.165 66.575 88.395 67.540 ;
        RECT 91.305 67.465 91.565 67.785 ;
        RECT 92.095 67.465 92.355 67.785 ;
        RECT 92.685 67.465 92.945 67.785 ;
        RECT 93.490 67.710 93.720 69.020 ;
        RECT 93.910 67.850 94.170 69.225 ;
        RECT 94.330 67.710 94.500 69.650 ;
        RECT 94.645 69.140 95.000 69.650 ;
        RECT 94.640 68.350 95.000 69.140 ;
        RECT 93.490 67.540 94.500 67.710 ;
        RECT 94.645 67.540 95.000 68.350 ;
        RECT 95.380 69.925 95.735 72.120 ;
        RECT 96.655 72.055 96.885 73.020 ;
        RECT 97.445 72.145 97.675 73.020 ;
        RECT 98.035 72.145 98.265 73.020 ;
        RECT 98.825 72.145 99.055 73.020 ;
        RECT 95.875 71.885 96.885 72.055 ;
        RECT 95.875 69.925 96.045 71.885 ;
        RECT 96.655 70.575 96.885 71.885 ;
        RECT 97.430 71.825 97.690 72.145 ;
        RECT 98.020 71.825 98.280 72.145 ;
        RECT 98.810 71.825 99.070 72.145 ;
        RECT 97.445 70.575 97.675 71.825 ;
        RECT 98.035 70.575 98.265 71.825 ;
        RECT 98.825 70.575 99.055 71.825 ;
        RECT 99.980 69.925 100.335 72.115 ;
        RECT 95.380 69.650 96.045 69.925 ;
        RECT 99.665 69.650 100.335 69.925 ;
        RECT 95.380 67.545 95.735 69.650 ;
        RECT 96.155 69.225 97.395 69.455 ;
        RECT 98.315 69.225 99.505 69.455 ;
        RECT 96.155 68.800 96.415 69.225 ;
        RECT 97.445 67.785 97.675 69.020 ;
        RECT 98.035 67.785 98.265 69.020 ;
        RECT 88.635 66.415 88.895 67.205 ;
        RECT 85.495 66.185 86.735 66.415 ;
        RECT 87.655 66.185 88.895 66.415 ;
        RECT 90.820 66.415 91.080 67.295 ;
        RECT 91.320 66.575 91.550 67.465 ;
        RECT 92.110 66.575 92.340 67.465 ;
        RECT 92.700 66.575 92.930 67.465 ;
        RECT 93.490 66.575 93.720 67.540 ;
        RECT 97.430 67.465 97.690 67.785 ;
        RECT 98.020 67.465 98.280 67.785 ;
        RECT 98.825 67.710 99.055 69.020 ;
        RECT 99.245 67.850 99.505 69.225 ;
        RECT 99.665 67.710 99.835 69.650 ;
        RECT 99.980 69.140 100.335 69.650 ;
        RECT 99.975 68.350 100.335 69.140 ;
        RECT 98.825 67.540 99.835 67.710 ;
        RECT 99.980 67.540 100.335 68.350 ;
        RECT 100.705 69.925 101.060 72.120 ;
        RECT 101.980 72.055 102.210 73.020 ;
        RECT 102.770 72.145 103.000 73.020 ;
        RECT 103.360 72.145 103.590 73.020 ;
        RECT 104.150 72.145 104.380 73.020 ;
        RECT 101.200 71.885 102.210 72.055 ;
        RECT 101.200 69.925 101.370 71.885 ;
        RECT 101.980 70.575 102.210 71.885 ;
        RECT 102.755 71.825 103.015 72.145 ;
        RECT 103.345 71.825 103.605 72.145 ;
        RECT 104.135 71.825 104.395 72.145 ;
        RECT 102.770 70.575 103.000 71.825 ;
        RECT 103.360 70.575 103.590 71.825 ;
        RECT 104.150 70.575 104.380 71.825 ;
        RECT 105.305 69.925 105.660 72.115 ;
        RECT 100.705 69.650 101.370 69.925 ;
        RECT 104.990 69.650 105.660 69.925 ;
        RECT 100.705 67.545 101.060 69.650 ;
        RECT 101.480 69.225 102.720 69.455 ;
        RECT 103.640 69.225 104.830 69.455 ;
        RECT 101.480 68.800 101.740 69.225 ;
        RECT 101.980 67.785 102.210 69.020 ;
        RECT 102.770 67.785 103.000 69.020 ;
        RECT 103.360 67.785 103.590 69.020 ;
        RECT 93.960 66.415 94.220 67.205 ;
        RECT 90.820 66.185 92.060 66.415 ;
        RECT 92.980 66.185 94.220 66.415 ;
        RECT 96.155 66.415 96.415 67.295 ;
        RECT 97.445 66.575 97.675 67.465 ;
        RECT 98.035 66.575 98.265 67.465 ;
        RECT 98.825 66.575 99.055 67.540 ;
        RECT 101.965 67.465 102.225 67.785 ;
        RECT 102.755 67.465 103.015 67.785 ;
        RECT 103.345 67.465 103.605 67.785 ;
        RECT 104.150 67.710 104.380 69.020 ;
        RECT 104.570 67.850 104.830 69.225 ;
        RECT 104.990 67.710 105.160 69.650 ;
        RECT 105.305 69.140 105.660 69.650 ;
        RECT 105.300 68.350 105.660 69.140 ;
        RECT 104.150 67.540 105.160 67.710 ;
        RECT 105.305 67.540 105.660 68.350 ;
        RECT 106.040 69.925 106.395 72.120 ;
        RECT 107.315 72.055 107.545 73.020 ;
        RECT 108.105 72.145 108.335 73.020 ;
        RECT 108.695 72.145 108.925 73.020 ;
        RECT 109.485 72.145 109.715 73.020 ;
        RECT 106.535 71.885 107.545 72.055 ;
        RECT 106.535 69.925 106.705 71.885 ;
        RECT 107.315 70.575 107.545 71.885 ;
        RECT 108.090 71.825 108.350 72.145 ;
        RECT 108.680 71.825 108.940 72.145 ;
        RECT 109.470 71.825 109.730 72.145 ;
        RECT 108.105 70.575 108.335 71.825 ;
        RECT 108.695 70.575 108.925 71.825 ;
        RECT 109.485 70.575 109.715 71.825 ;
        RECT 110.640 69.925 110.995 72.115 ;
        RECT 106.040 69.650 106.705 69.925 ;
        RECT 110.325 69.650 110.995 69.925 ;
        RECT 106.040 67.545 106.395 69.650 ;
        RECT 106.815 69.225 108.055 69.455 ;
        RECT 108.975 69.225 110.165 69.455 ;
        RECT 106.815 68.800 107.075 69.225 ;
        RECT 107.315 67.785 107.545 69.020 ;
        RECT 108.105 67.785 108.335 69.020 ;
        RECT 108.695 67.785 108.925 69.020 ;
        RECT 99.295 66.415 99.555 67.205 ;
        RECT 96.155 66.185 97.395 66.415 ;
        RECT 98.315 66.185 99.555 66.415 ;
        RECT 101.480 66.415 101.740 67.295 ;
        RECT 101.980 66.575 102.210 67.465 ;
        RECT 102.770 66.575 103.000 67.465 ;
        RECT 103.360 66.575 103.590 67.465 ;
        RECT 104.150 66.575 104.380 67.540 ;
        RECT 107.300 67.465 107.560 67.785 ;
        RECT 108.090 67.465 108.350 67.785 ;
        RECT 108.680 67.465 108.940 67.785 ;
        RECT 109.485 67.710 109.715 69.020 ;
        RECT 109.905 67.850 110.165 69.225 ;
        RECT 110.325 67.710 110.495 69.650 ;
        RECT 110.640 69.140 110.995 69.650 ;
        RECT 110.635 68.350 110.995 69.140 ;
        RECT 109.485 67.540 110.495 67.710 ;
        RECT 110.640 67.540 110.995 68.350 ;
        RECT 111.365 69.925 111.720 72.120 ;
        RECT 112.640 72.055 112.870 73.020 ;
        RECT 113.430 72.145 113.660 73.020 ;
        RECT 114.020 72.145 114.250 73.020 ;
        RECT 114.810 72.145 115.040 73.020 ;
        RECT 111.860 71.885 112.870 72.055 ;
        RECT 111.860 69.925 112.030 71.885 ;
        RECT 112.640 70.575 112.870 71.885 ;
        RECT 113.415 71.825 113.675 72.145 ;
        RECT 114.005 71.825 114.265 72.145 ;
        RECT 114.795 71.825 115.055 72.145 ;
        RECT 113.430 70.575 113.660 71.825 ;
        RECT 114.020 70.575 114.250 71.825 ;
        RECT 114.810 70.575 115.040 71.825 ;
        RECT 115.965 69.925 116.320 72.115 ;
        RECT 111.365 69.650 112.030 69.925 ;
        RECT 115.650 69.650 116.320 69.925 ;
        RECT 111.365 67.545 111.720 69.650 ;
        RECT 112.140 69.225 113.380 69.455 ;
        RECT 114.300 69.225 115.490 69.455 ;
        RECT 112.140 68.800 112.400 69.225 ;
        RECT 112.640 67.785 112.870 69.020 ;
        RECT 113.430 67.785 113.660 69.020 ;
        RECT 114.020 67.785 114.250 69.020 ;
        RECT 104.620 66.415 104.880 67.205 ;
        RECT 101.480 66.185 102.720 66.415 ;
        RECT 103.640 66.185 104.880 66.415 ;
        RECT 106.815 66.415 107.075 67.295 ;
        RECT 107.315 66.575 107.545 67.465 ;
        RECT 108.105 66.575 108.335 67.465 ;
        RECT 108.695 66.575 108.925 67.465 ;
        RECT 109.485 66.575 109.715 67.540 ;
        RECT 112.625 67.465 112.885 67.785 ;
        RECT 113.415 67.465 113.675 67.785 ;
        RECT 114.005 67.465 114.265 67.785 ;
        RECT 114.810 67.710 115.040 69.020 ;
        RECT 115.230 67.850 115.490 69.225 ;
        RECT 115.650 67.710 115.820 69.650 ;
        RECT 115.965 69.140 116.320 69.650 ;
        RECT 115.960 68.350 116.320 69.140 ;
        RECT 114.810 67.540 115.820 67.710 ;
        RECT 115.965 67.540 116.320 68.350 ;
        RECT 116.700 69.925 117.055 72.120 ;
        RECT 117.975 72.055 118.205 73.020 ;
        RECT 118.765 72.145 118.995 73.020 ;
        RECT 119.355 72.145 119.585 73.020 ;
        RECT 120.145 72.145 120.375 73.020 ;
        RECT 117.195 71.885 118.205 72.055 ;
        RECT 117.195 69.925 117.365 71.885 ;
        RECT 117.975 70.575 118.205 71.885 ;
        RECT 118.750 71.825 119.010 72.145 ;
        RECT 119.340 71.825 119.600 72.145 ;
        RECT 120.130 71.825 120.390 72.145 ;
        RECT 118.765 70.575 118.995 71.825 ;
        RECT 119.355 70.575 119.585 71.825 ;
        RECT 120.145 70.575 120.375 71.825 ;
        RECT 121.300 69.925 121.655 72.115 ;
        RECT 116.700 69.650 117.365 69.925 ;
        RECT 120.985 69.650 121.655 69.925 ;
        RECT 116.700 67.545 117.055 69.650 ;
        RECT 119.635 69.225 120.825 69.455 ;
        RECT 117.975 67.785 118.205 69.020 ;
        RECT 118.765 67.785 118.995 69.020 ;
        RECT 119.355 67.785 119.585 69.020 ;
        RECT 109.955 66.415 110.215 67.205 ;
        RECT 106.815 66.185 108.055 66.415 ;
        RECT 108.975 66.185 110.215 66.415 ;
        RECT 112.140 66.415 112.400 67.295 ;
        RECT 112.640 66.575 112.870 67.465 ;
        RECT 113.430 66.575 113.660 67.465 ;
        RECT 114.020 66.575 114.250 67.465 ;
        RECT 114.810 66.575 115.040 67.540 ;
        RECT 117.960 67.465 118.220 67.785 ;
        RECT 118.750 67.465 119.010 67.785 ;
        RECT 119.340 67.465 119.600 67.785 ;
        RECT 120.145 67.710 120.375 69.020 ;
        RECT 120.565 67.850 120.825 69.225 ;
        RECT 120.985 67.710 121.155 69.650 ;
        RECT 121.300 69.140 121.655 69.650 ;
        RECT 121.295 68.350 121.655 69.140 ;
        RECT 120.145 67.540 121.155 67.710 ;
        RECT 121.300 67.540 121.655 68.350 ;
        RECT 122.025 69.925 122.380 72.135 ;
        RECT 123.300 72.055 123.530 73.020 ;
        RECT 124.090 72.145 124.320 73.020 ;
        RECT 124.680 72.145 124.910 73.020 ;
        RECT 125.470 72.145 125.700 73.020 ;
        RECT 122.520 71.885 123.530 72.055 ;
        RECT 122.520 69.925 122.690 71.885 ;
        RECT 123.300 70.575 123.530 71.885 ;
        RECT 124.075 71.825 124.335 72.145 ;
        RECT 124.665 71.825 124.925 72.145 ;
        RECT 125.455 71.825 125.715 72.145 ;
        RECT 124.090 70.575 124.320 71.825 ;
        RECT 124.680 70.575 124.910 71.825 ;
        RECT 125.470 70.575 125.700 71.825 ;
        RECT 126.625 69.925 126.980 72.135 ;
        RECT 122.025 69.650 122.690 69.925 ;
        RECT 126.310 69.650 126.980 69.925 ;
        RECT 122.025 67.560 122.380 69.650 ;
        RECT 123.300 67.785 123.530 69.020 ;
        RECT 124.090 67.785 124.320 69.020 ;
        RECT 124.680 67.785 124.910 69.020 ;
        RECT 122.115 67.540 122.375 67.560 ;
        RECT 115.280 66.415 115.540 67.205 ;
        RECT 117.975 66.575 118.205 67.465 ;
        RECT 118.765 66.575 118.995 67.465 ;
        RECT 119.355 66.575 119.585 67.465 ;
        RECT 120.145 66.575 120.375 67.540 ;
        RECT 123.285 67.465 123.545 67.785 ;
        RECT 124.075 67.465 124.335 67.785 ;
        RECT 124.665 67.465 124.925 67.785 ;
        RECT 125.470 67.710 125.700 69.020 ;
        RECT 126.310 67.710 126.480 69.650 ;
        RECT 126.625 67.855 126.980 69.650 ;
        RECT 125.470 67.540 126.480 67.710 ;
        RECT 126.620 67.560 126.980 67.855 ;
        RECT 120.615 66.415 120.875 67.205 ;
        RECT 123.300 66.575 123.530 67.465 ;
        RECT 124.090 66.575 124.320 67.465 ;
        RECT 124.680 66.575 124.910 67.465 ;
        RECT 125.470 66.575 125.700 67.540 ;
        RECT 126.620 67.535 126.880 67.560 ;
        RECT 112.140 66.185 113.380 66.415 ;
        RECT 114.300 66.185 115.540 66.415 ;
        RECT 119.635 66.185 120.875 66.415 ;
        RECT 22.725 65.675 22.985 65.680 ;
        RECT 10.510 64.155 10.810 65.605 ;
        RECT 15.985 65.440 23.050 65.675 ;
        RECT 37.520 65.645 38.760 65.875 ;
        RECT 39.680 65.645 40.920 65.875 ;
        RECT 11.745 65.055 13.345 65.345 ;
        RECT 14.165 65.055 20.945 65.290 ;
        RECT 16.040 64.870 17.645 64.900 ;
        RECT 21.425 64.870 23.050 65.440 ;
        RECT 15.985 64.635 23.050 64.870 ;
        RECT 16.040 64.610 17.645 64.635 ;
        RECT 31.420 62.390 31.775 64.600 ;
        RECT 32.695 64.520 32.925 65.485 ;
        RECT 33.485 64.610 33.715 65.485 ;
        RECT 34.075 64.610 34.305 65.485 ;
        RECT 34.865 64.610 35.095 65.485 ;
        RECT 37.520 64.950 37.780 65.645 ;
        RECT 31.915 64.350 32.925 64.520 ;
        RECT 31.915 62.390 32.085 64.350 ;
        RECT 32.695 63.040 32.925 64.350 ;
        RECT 33.470 64.290 33.730 64.610 ;
        RECT 34.060 64.290 34.320 64.610 ;
        RECT 34.850 64.290 35.110 64.610 ;
        RECT 33.485 63.040 33.715 64.290 ;
        RECT 34.075 63.040 34.305 64.290 ;
        RECT 34.865 63.040 35.095 64.290 ;
        RECT 36.020 62.390 36.375 64.600 ;
        RECT 31.420 62.115 32.085 62.390 ;
        RECT 35.705 62.115 36.375 62.390 ;
        RECT 10.500 60.610 10.820 61.095 ;
        RECT 16.115 60.720 23.440 60.955 ;
        RECT 10.500 60.280 11.960 60.610 ;
        RECT 10.500 60.060 10.820 60.280 ;
        RECT 12.400 59.535 12.720 60.525 ;
        RECT 14.585 60.280 16.005 60.605 ;
        RECT 19.990 60.150 23.440 60.720 ;
        RECT 16.115 59.915 23.440 60.150 ;
        RECT 31.420 60.025 31.775 62.115 ;
        RECT 32.695 60.250 32.925 61.485 ;
        RECT 33.485 60.250 33.715 61.485 ;
        RECT 34.075 60.250 34.305 61.485 ;
        RECT 32.680 59.930 32.940 60.250 ;
        RECT 33.470 59.930 33.730 60.250 ;
        RECT 34.060 59.930 34.320 60.250 ;
        RECT 34.865 60.175 35.095 61.485 ;
        RECT 35.705 60.175 35.875 62.115 ;
        RECT 34.865 60.005 35.875 60.175 ;
        RECT 36.020 60.025 36.375 62.115 ;
        RECT 36.745 62.390 37.100 64.585 ;
        RECT 38.020 64.520 38.250 65.485 ;
        RECT 38.810 64.610 39.040 65.485 ;
        RECT 39.400 64.610 39.630 65.485 ;
        RECT 40.190 64.610 40.420 65.485 ;
        RECT 40.660 64.855 40.920 65.645 ;
        RECT 42.855 65.645 44.095 65.875 ;
        RECT 45.015 65.645 46.255 65.875 ;
        RECT 42.855 64.950 43.115 65.645 ;
        RECT 37.240 64.350 38.250 64.520 ;
        RECT 37.240 62.390 37.410 64.350 ;
        RECT 37.570 62.835 37.830 63.970 ;
        RECT 38.020 63.040 38.250 64.350 ;
        RECT 38.795 64.290 39.055 64.610 ;
        RECT 39.385 64.290 39.645 64.610 ;
        RECT 40.175 64.290 40.435 64.610 ;
        RECT 38.810 63.040 39.040 64.290 ;
        RECT 39.400 63.040 39.630 64.290 ;
        RECT 40.190 63.040 40.420 64.290 ;
        RECT 40.660 62.835 40.920 63.340 ;
        RECT 37.570 62.605 38.760 62.835 ;
        RECT 39.680 62.605 40.920 62.835 ;
        RECT 41.345 62.390 41.700 64.580 ;
        RECT 36.745 62.115 37.410 62.390 ;
        RECT 41.030 62.115 41.700 62.390 ;
        RECT 36.745 60.010 37.100 62.115 ;
        RECT 37.520 61.690 38.760 61.920 ;
        RECT 39.680 61.690 40.870 61.920 ;
        RECT 37.520 61.265 37.780 61.690 ;
        RECT 38.020 60.250 38.250 61.485 ;
        RECT 38.810 60.250 39.040 61.485 ;
        RECT 39.400 60.250 39.630 61.485 ;
        RECT 12.425 59.520 12.715 59.535 ;
        RECT 32.695 59.040 32.925 59.930 ;
        RECT 33.485 59.040 33.715 59.930 ;
        RECT 34.075 59.040 34.305 59.930 ;
        RECT 34.865 59.040 35.095 60.005 ;
        RECT 38.005 59.930 38.265 60.250 ;
        RECT 38.795 59.930 39.055 60.250 ;
        RECT 39.385 59.930 39.645 60.250 ;
        RECT 40.190 60.175 40.420 61.485 ;
        RECT 40.610 60.615 40.870 61.690 ;
        RECT 41.030 60.175 41.200 62.115 ;
        RECT 40.190 60.005 41.200 60.175 ;
        RECT 41.345 60.005 41.700 62.115 ;
        RECT 42.080 62.390 42.435 64.585 ;
        RECT 43.355 64.520 43.585 65.485 ;
        RECT 44.145 64.610 44.375 65.485 ;
        RECT 44.735 64.610 44.965 65.485 ;
        RECT 45.525 64.610 45.755 65.485 ;
        RECT 45.995 64.855 46.255 65.645 ;
        RECT 48.180 65.645 49.420 65.875 ;
        RECT 50.340 65.645 51.580 65.875 ;
        RECT 48.180 64.950 48.440 65.645 ;
        RECT 42.575 64.350 43.585 64.520 ;
        RECT 42.575 62.390 42.745 64.350 ;
        RECT 42.905 62.835 43.165 63.970 ;
        RECT 43.355 63.040 43.585 64.350 ;
        RECT 44.130 64.290 44.390 64.610 ;
        RECT 44.720 64.290 44.980 64.610 ;
        RECT 45.510 64.290 45.770 64.610 ;
        RECT 44.145 63.040 44.375 64.290 ;
        RECT 44.735 63.040 44.965 64.290 ;
        RECT 45.525 63.040 45.755 64.290 ;
        RECT 45.995 62.835 46.255 63.340 ;
        RECT 42.905 62.605 44.095 62.835 ;
        RECT 45.015 62.605 46.255 62.835 ;
        RECT 46.680 62.390 47.035 64.580 ;
        RECT 42.080 62.115 42.745 62.390 ;
        RECT 46.365 62.115 47.035 62.390 ;
        RECT 42.080 60.010 42.435 62.115 ;
        RECT 42.855 61.690 44.095 61.920 ;
        RECT 45.015 61.690 46.205 61.920 ;
        RECT 42.855 61.265 43.115 61.690 ;
        RECT 43.355 60.250 43.585 61.485 ;
        RECT 44.145 60.250 44.375 61.485 ;
        RECT 44.735 60.250 44.965 61.485 ;
        RECT 37.520 58.880 37.780 59.760 ;
        RECT 38.020 59.040 38.250 59.930 ;
        RECT 38.810 59.040 39.040 59.930 ;
        RECT 39.400 59.040 39.630 59.930 ;
        RECT 40.190 59.040 40.420 60.005 ;
        RECT 43.340 59.930 43.600 60.250 ;
        RECT 44.130 59.930 44.390 60.250 ;
        RECT 44.720 59.930 44.980 60.250 ;
        RECT 45.525 60.175 45.755 61.485 ;
        RECT 45.945 60.615 46.205 61.690 ;
        RECT 46.365 60.175 46.535 62.115 ;
        RECT 45.525 60.005 46.535 60.175 ;
        RECT 46.680 60.005 47.035 62.115 ;
        RECT 47.405 62.390 47.760 64.585 ;
        RECT 48.680 64.520 48.910 65.485 ;
        RECT 49.470 64.610 49.700 65.485 ;
        RECT 50.060 64.610 50.290 65.485 ;
        RECT 50.850 64.610 51.080 65.485 ;
        RECT 51.320 64.855 51.580 65.645 ;
        RECT 53.515 65.645 54.755 65.875 ;
        RECT 55.675 65.645 56.915 65.875 ;
        RECT 53.515 64.950 53.775 65.645 ;
        RECT 47.900 64.350 48.910 64.520 ;
        RECT 47.900 62.390 48.070 64.350 ;
        RECT 48.230 62.835 48.490 63.970 ;
        RECT 48.680 63.040 48.910 64.350 ;
        RECT 49.455 64.290 49.715 64.610 ;
        RECT 50.045 64.290 50.305 64.610 ;
        RECT 50.835 64.290 51.095 64.610 ;
        RECT 49.470 63.040 49.700 64.290 ;
        RECT 50.060 63.040 50.290 64.290 ;
        RECT 50.850 63.040 51.080 64.290 ;
        RECT 51.320 62.835 51.580 63.340 ;
        RECT 48.230 62.605 49.420 62.835 ;
        RECT 50.340 62.605 51.580 62.835 ;
        RECT 52.005 62.390 52.360 64.580 ;
        RECT 47.405 62.115 48.070 62.390 ;
        RECT 51.690 62.115 52.360 62.390 ;
        RECT 47.405 60.010 47.760 62.115 ;
        RECT 48.180 61.690 49.420 61.920 ;
        RECT 50.340 61.690 51.530 61.920 ;
        RECT 48.180 61.265 48.440 61.690 ;
        RECT 48.680 60.250 48.910 61.485 ;
        RECT 49.470 60.250 49.700 61.485 ;
        RECT 50.060 60.250 50.290 61.485 ;
        RECT 40.660 58.880 40.920 59.670 ;
        RECT 37.520 58.650 38.760 58.880 ;
        RECT 39.680 58.650 40.920 58.880 ;
        RECT 42.855 58.880 43.115 59.760 ;
        RECT 43.355 59.040 43.585 59.930 ;
        RECT 44.145 59.040 44.375 59.930 ;
        RECT 44.735 59.040 44.965 59.930 ;
        RECT 45.525 59.040 45.755 60.005 ;
        RECT 48.665 59.930 48.925 60.250 ;
        RECT 49.455 59.930 49.715 60.250 ;
        RECT 50.045 59.930 50.305 60.250 ;
        RECT 50.850 60.175 51.080 61.485 ;
        RECT 51.270 60.615 51.530 61.690 ;
        RECT 51.690 60.175 51.860 62.115 ;
        RECT 50.850 60.005 51.860 60.175 ;
        RECT 52.005 60.005 52.360 62.115 ;
        RECT 52.740 62.390 53.095 64.585 ;
        RECT 54.015 64.520 54.245 65.485 ;
        RECT 54.805 64.610 55.035 65.485 ;
        RECT 55.395 64.610 55.625 65.485 ;
        RECT 56.185 64.610 56.415 65.485 ;
        RECT 56.655 64.855 56.915 65.645 ;
        RECT 58.840 65.645 60.080 65.875 ;
        RECT 61.000 65.645 62.240 65.875 ;
        RECT 58.840 64.950 59.100 65.645 ;
        RECT 53.235 64.350 54.245 64.520 ;
        RECT 53.235 62.390 53.405 64.350 ;
        RECT 53.565 62.835 53.825 63.970 ;
        RECT 54.015 63.040 54.245 64.350 ;
        RECT 54.790 64.290 55.050 64.610 ;
        RECT 55.380 64.290 55.640 64.610 ;
        RECT 56.170 64.290 56.430 64.610 ;
        RECT 54.805 63.040 55.035 64.290 ;
        RECT 55.395 63.040 55.625 64.290 ;
        RECT 56.185 63.040 56.415 64.290 ;
        RECT 56.655 62.835 56.915 63.340 ;
        RECT 53.565 62.605 54.755 62.835 ;
        RECT 55.675 62.605 56.915 62.835 ;
        RECT 57.340 62.390 57.695 64.580 ;
        RECT 52.740 62.115 53.405 62.390 ;
        RECT 57.025 62.115 57.695 62.390 ;
        RECT 52.740 60.010 53.095 62.115 ;
        RECT 53.515 61.690 54.755 61.920 ;
        RECT 55.675 61.690 56.865 61.920 ;
        RECT 53.515 61.265 53.775 61.690 ;
        RECT 54.015 60.250 54.245 61.485 ;
        RECT 54.805 60.250 55.035 61.485 ;
        RECT 55.395 60.250 55.625 61.485 ;
        RECT 45.995 58.880 46.255 59.670 ;
        RECT 42.855 58.650 44.095 58.880 ;
        RECT 45.015 58.650 46.255 58.880 ;
        RECT 48.180 58.880 48.440 59.760 ;
        RECT 48.680 59.040 48.910 59.930 ;
        RECT 49.470 59.040 49.700 59.930 ;
        RECT 50.060 59.040 50.290 59.930 ;
        RECT 50.850 59.040 51.080 60.005 ;
        RECT 54.000 59.930 54.260 60.250 ;
        RECT 54.790 59.930 55.050 60.250 ;
        RECT 55.380 59.930 55.640 60.250 ;
        RECT 56.185 60.175 56.415 61.485 ;
        RECT 56.605 60.615 56.865 61.690 ;
        RECT 57.025 60.175 57.195 62.115 ;
        RECT 56.185 60.005 57.195 60.175 ;
        RECT 57.340 60.005 57.695 62.115 ;
        RECT 58.065 62.390 58.420 64.585 ;
        RECT 59.340 64.520 59.570 65.485 ;
        RECT 60.130 64.610 60.360 65.485 ;
        RECT 60.720 64.610 60.950 65.485 ;
        RECT 61.510 64.610 61.740 65.485 ;
        RECT 61.980 64.855 62.240 65.645 ;
        RECT 64.175 65.645 65.415 65.875 ;
        RECT 66.335 65.645 67.575 65.875 ;
        RECT 64.175 64.950 64.435 65.645 ;
        RECT 58.560 64.350 59.570 64.520 ;
        RECT 58.560 62.390 58.730 64.350 ;
        RECT 58.890 62.835 59.150 63.970 ;
        RECT 59.340 63.040 59.570 64.350 ;
        RECT 60.115 64.290 60.375 64.610 ;
        RECT 60.705 64.290 60.965 64.610 ;
        RECT 61.495 64.290 61.755 64.610 ;
        RECT 60.130 63.040 60.360 64.290 ;
        RECT 60.720 63.040 60.950 64.290 ;
        RECT 61.510 63.040 61.740 64.290 ;
        RECT 61.980 62.835 62.240 63.340 ;
        RECT 58.890 62.605 60.080 62.835 ;
        RECT 61.000 62.605 62.240 62.835 ;
        RECT 62.665 62.390 63.020 64.580 ;
        RECT 58.065 62.115 58.730 62.390 ;
        RECT 62.350 62.115 63.020 62.390 ;
        RECT 58.065 60.010 58.420 62.115 ;
        RECT 58.840 61.690 60.080 61.920 ;
        RECT 61.000 61.690 62.190 61.920 ;
        RECT 58.840 61.265 59.100 61.690 ;
        RECT 59.340 60.250 59.570 61.485 ;
        RECT 60.130 60.250 60.360 61.485 ;
        RECT 60.720 60.250 60.950 61.485 ;
        RECT 51.320 58.880 51.580 59.670 ;
        RECT 48.180 58.650 49.420 58.880 ;
        RECT 50.340 58.650 51.580 58.880 ;
        RECT 53.515 58.880 53.775 59.760 ;
        RECT 54.015 59.040 54.245 59.930 ;
        RECT 54.805 59.040 55.035 59.930 ;
        RECT 55.395 59.040 55.625 59.930 ;
        RECT 56.185 59.040 56.415 60.005 ;
        RECT 59.325 59.930 59.585 60.250 ;
        RECT 60.115 59.930 60.375 60.250 ;
        RECT 60.705 59.930 60.965 60.250 ;
        RECT 61.510 60.175 61.740 61.485 ;
        RECT 61.930 60.615 62.190 61.690 ;
        RECT 62.350 60.175 62.520 62.115 ;
        RECT 61.510 60.005 62.520 60.175 ;
        RECT 62.665 60.005 63.020 62.115 ;
        RECT 63.400 62.390 63.755 64.585 ;
        RECT 64.675 64.520 64.905 65.485 ;
        RECT 65.465 64.610 65.695 65.485 ;
        RECT 66.055 64.610 66.285 65.485 ;
        RECT 66.845 64.610 67.075 65.485 ;
        RECT 67.315 64.855 67.575 65.645 ;
        RECT 69.500 65.645 70.740 65.875 ;
        RECT 71.660 65.645 72.900 65.875 ;
        RECT 69.500 64.950 69.760 65.645 ;
        RECT 63.895 64.350 64.905 64.520 ;
        RECT 63.895 62.390 64.065 64.350 ;
        RECT 64.225 62.835 64.485 63.970 ;
        RECT 64.675 63.040 64.905 64.350 ;
        RECT 65.450 64.290 65.710 64.610 ;
        RECT 66.040 64.290 66.300 64.610 ;
        RECT 66.830 64.290 67.090 64.610 ;
        RECT 65.465 63.040 65.695 64.290 ;
        RECT 66.055 63.040 66.285 64.290 ;
        RECT 66.845 63.040 67.075 64.290 ;
        RECT 67.315 62.835 67.575 63.340 ;
        RECT 64.225 62.605 65.415 62.835 ;
        RECT 66.335 62.605 67.575 62.835 ;
        RECT 68.000 62.390 68.355 64.580 ;
        RECT 63.400 62.115 64.065 62.390 ;
        RECT 67.685 62.115 68.355 62.390 ;
        RECT 63.400 60.010 63.755 62.115 ;
        RECT 64.175 61.690 65.415 61.920 ;
        RECT 66.335 61.690 67.525 61.920 ;
        RECT 64.175 61.265 64.435 61.690 ;
        RECT 64.675 60.250 64.905 61.485 ;
        RECT 65.465 60.250 65.695 61.485 ;
        RECT 66.055 60.250 66.285 61.485 ;
        RECT 56.655 58.880 56.915 59.670 ;
        RECT 53.515 58.650 54.755 58.880 ;
        RECT 55.675 58.650 56.915 58.880 ;
        RECT 58.840 58.880 59.100 59.760 ;
        RECT 59.340 59.040 59.570 59.930 ;
        RECT 60.130 59.040 60.360 59.930 ;
        RECT 60.720 59.040 60.950 59.930 ;
        RECT 61.510 59.040 61.740 60.005 ;
        RECT 64.660 59.930 64.920 60.250 ;
        RECT 65.450 59.930 65.710 60.250 ;
        RECT 66.040 59.930 66.300 60.250 ;
        RECT 66.845 60.175 67.075 61.485 ;
        RECT 67.265 60.615 67.525 61.690 ;
        RECT 67.685 60.175 67.855 62.115 ;
        RECT 66.845 60.005 67.855 60.175 ;
        RECT 68.000 60.005 68.355 62.115 ;
        RECT 68.725 62.390 69.080 64.585 ;
        RECT 70.000 64.520 70.230 65.485 ;
        RECT 70.790 64.610 71.020 65.485 ;
        RECT 71.380 64.610 71.610 65.485 ;
        RECT 72.170 64.610 72.400 65.485 ;
        RECT 72.640 64.855 72.900 65.645 ;
        RECT 74.835 65.645 76.075 65.875 ;
        RECT 76.995 65.645 78.235 65.875 ;
        RECT 74.835 64.950 75.095 65.645 ;
        RECT 69.220 64.350 70.230 64.520 ;
        RECT 69.220 62.390 69.390 64.350 ;
        RECT 69.550 62.835 69.810 63.970 ;
        RECT 70.000 63.040 70.230 64.350 ;
        RECT 70.775 64.290 71.035 64.610 ;
        RECT 71.365 64.290 71.625 64.610 ;
        RECT 72.155 64.290 72.415 64.610 ;
        RECT 70.790 63.040 71.020 64.290 ;
        RECT 71.380 63.040 71.610 64.290 ;
        RECT 72.170 63.040 72.400 64.290 ;
        RECT 72.640 62.835 72.900 63.340 ;
        RECT 69.550 62.605 70.740 62.835 ;
        RECT 71.660 62.605 72.900 62.835 ;
        RECT 73.325 62.390 73.680 64.580 ;
        RECT 68.725 62.115 69.390 62.390 ;
        RECT 73.010 62.115 73.680 62.390 ;
        RECT 68.725 60.010 69.080 62.115 ;
        RECT 69.500 61.690 70.740 61.920 ;
        RECT 71.660 61.690 72.850 61.920 ;
        RECT 69.500 61.265 69.760 61.690 ;
        RECT 70.000 60.250 70.230 61.485 ;
        RECT 70.790 60.250 71.020 61.485 ;
        RECT 71.380 60.250 71.610 61.485 ;
        RECT 61.980 58.880 62.240 59.670 ;
        RECT 58.840 58.650 60.080 58.880 ;
        RECT 61.000 58.650 62.240 58.880 ;
        RECT 64.175 58.880 64.435 59.760 ;
        RECT 64.675 59.040 64.905 59.930 ;
        RECT 65.465 59.040 65.695 59.930 ;
        RECT 66.055 59.040 66.285 59.930 ;
        RECT 66.845 59.040 67.075 60.005 ;
        RECT 69.985 59.930 70.245 60.250 ;
        RECT 70.775 59.930 71.035 60.250 ;
        RECT 71.365 59.930 71.625 60.250 ;
        RECT 72.170 60.175 72.400 61.485 ;
        RECT 72.590 60.615 72.850 61.690 ;
        RECT 73.010 60.175 73.180 62.115 ;
        RECT 72.170 60.005 73.180 60.175 ;
        RECT 73.325 60.005 73.680 62.115 ;
        RECT 74.060 62.390 74.415 64.585 ;
        RECT 75.335 64.520 75.565 65.485 ;
        RECT 76.125 64.610 76.355 65.485 ;
        RECT 76.715 64.610 76.945 65.485 ;
        RECT 77.505 64.610 77.735 65.485 ;
        RECT 77.975 64.855 78.235 65.645 ;
        RECT 80.160 65.645 81.400 65.875 ;
        RECT 82.320 65.645 83.560 65.875 ;
        RECT 80.160 64.950 80.420 65.645 ;
        RECT 74.555 64.350 75.565 64.520 ;
        RECT 74.555 62.390 74.725 64.350 ;
        RECT 74.885 62.835 75.145 63.970 ;
        RECT 75.335 63.040 75.565 64.350 ;
        RECT 76.110 64.290 76.370 64.610 ;
        RECT 76.700 64.290 76.960 64.610 ;
        RECT 77.490 64.290 77.750 64.610 ;
        RECT 76.125 63.040 76.355 64.290 ;
        RECT 76.715 63.040 76.945 64.290 ;
        RECT 77.505 63.040 77.735 64.290 ;
        RECT 77.975 62.835 78.235 63.340 ;
        RECT 74.885 62.605 76.075 62.835 ;
        RECT 76.995 62.605 78.235 62.835 ;
        RECT 78.660 62.390 79.015 64.580 ;
        RECT 74.060 62.115 74.725 62.390 ;
        RECT 78.345 62.115 79.015 62.390 ;
        RECT 74.060 60.010 74.415 62.115 ;
        RECT 74.835 61.690 76.075 61.920 ;
        RECT 76.995 61.690 78.185 61.920 ;
        RECT 74.835 61.265 75.095 61.690 ;
        RECT 75.335 60.250 75.565 61.485 ;
        RECT 76.125 60.250 76.355 61.485 ;
        RECT 76.715 60.250 76.945 61.485 ;
        RECT 67.315 58.880 67.575 59.670 ;
        RECT 64.175 58.650 65.415 58.880 ;
        RECT 66.335 58.650 67.575 58.880 ;
        RECT 69.500 58.880 69.760 59.760 ;
        RECT 70.000 59.040 70.230 59.930 ;
        RECT 70.790 59.040 71.020 59.930 ;
        RECT 71.380 59.040 71.610 59.930 ;
        RECT 72.170 59.040 72.400 60.005 ;
        RECT 75.320 59.930 75.580 60.250 ;
        RECT 76.110 59.930 76.370 60.250 ;
        RECT 76.700 59.930 76.960 60.250 ;
        RECT 77.505 60.175 77.735 61.485 ;
        RECT 77.925 60.615 78.185 61.690 ;
        RECT 78.345 60.175 78.515 62.115 ;
        RECT 77.505 60.005 78.515 60.175 ;
        RECT 78.660 60.005 79.015 62.115 ;
        RECT 79.385 62.390 79.740 64.585 ;
        RECT 80.660 64.520 80.890 65.485 ;
        RECT 81.450 64.610 81.680 65.485 ;
        RECT 82.040 64.610 82.270 65.485 ;
        RECT 82.830 64.610 83.060 65.485 ;
        RECT 83.300 64.855 83.560 65.645 ;
        RECT 85.495 65.645 86.735 65.875 ;
        RECT 87.655 65.645 88.895 65.875 ;
        RECT 85.495 64.950 85.755 65.645 ;
        RECT 79.880 64.350 80.890 64.520 ;
        RECT 79.880 62.390 80.050 64.350 ;
        RECT 80.210 62.835 80.470 63.970 ;
        RECT 80.660 63.040 80.890 64.350 ;
        RECT 81.435 64.290 81.695 64.610 ;
        RECT 82.025 64.290 82.285 64.610 ;
        RECT 82.815 64.290 83.075 64.610 ;
        RECT 81.450 63.040 81.680 64.290 ;
        RECT 82.040 63.040 82.270 64.290 ;
        RECT 82.830 63.040 83.060 64.290 ;
        RECT 83.300 62.835 83.560 63.340 ;
        RECT 80.210 62.605 81.400 62.835 ;
        RECT 82.320 62.605 83.560 62.835 ;
        RECT 83.985 62.390 84.340 64.580 ;
        RECT 79.385 62.115 80.050 62.390 ;
        RECT 83.670 62.115 84.340 62.390 ;
        RECT 79.385 60.010 79.740 62.115 ;
        RECT 80.160 61.690 81.400 61.920 ;
        RECT 82.320 61.690 83.510 61.920 ;
        RECT 80.160 61.265 80.420 61.690 ;
        RECT 80.660 60.250 80.890 61.485 ;
        RECT 81.450 60.250 81.680 61.485 ;
        RECT 82.040 60.250 82.270 61.485 ;
        RECT 72.640 58.880 72.900 59.670 ;
        RECT 69.500 58.650 70.740 58.880 ;
        RECT 71.660 58.650 72.900 58.880 ;
        RECT 74.835 58.880 75.095 59.760 ;
        RECT 75.335 59.040 75.565 59.930 ;
        RECT 76.125 59.040 76.355 59.930 ;
        RECT 76.715 59.040 76.945 59.930 ;
        RECT 77.505 59.040 77.735 60.005 ;
        RECT 80.645 59.930 80.905 60.250 ;
        RECT 81.435 59.930 81.695 60.250 ;
        RECT 82.025 59.930 82.285 60.250 ;
        RECT 82.830 60.175 83.060 61.485 ;
        RECT 83.250 60.615 83.510 61.690 ;
        RECT 83.670 60.175 83.840 62.115 ;
        RECT 82.830 60.005 83.840 60.175 ;
        RECT 83.985 60.005 84.340 62.115 ;
        RECT 84.720 62.390 85.075 64.585 ;
        RECT 85.995 64.520 86.225 65.485 ;
        RECT 86.785 64.610 87.015 65.485 ;
        RECT 87.375 64.610 87.605 65.485 ;
        RECT 88.165 64.610 88.395 65.485 ;
        RECT 88.635 64.855 88.895 65.645 ;
        RECT 90.820 65.645 92.060 65.875 ;
        RECT 92.980 65.645 94.220 65.875 ;
        RECT 90.820 64.950 91.080 65.645 ;
        RECT 85.215 64.350 86.225 64.520 ;
        RECT 85.215 62.390 85.385 64.350 ;
        RECT 85.545 62.835 85.805 63.970 ;
        RECT 85.995 63.040 86.225 64.350 ;
        RECT 86.770 64.290 87.030 64.610 ;
        RECT 87.360 64.290 87.620 64.610 ;
        RECT 88.150 64.290 88.410 64.610 ;
        RECT 86.785 63.040 87.015 64.290 ;
        RECT 87.375 63.040 87.605 64.290 ;
        RECT 88.165 63.040 88.395 64.290 ;
        RECT 88.635 62.835 88.895 63.340 ;
        RECT 85.545 62.605 86.735 62.835 ;
        RECT 87.655 62.605 88.895 62.835 ;
        RECT 89.320 62.390 89.675 64.580 ;
        RECT 84.720 62.115 85.385 62.390 ;
        RECT 89.005 62.115 89.675 62.390 ;
        RECT 84.720 60.010 85.075 62.115 ;
        RECT 85.495 61.690 86.735 61.920 ;
        RECT 87.655 61.690 88.845 61.920 ;
        RECT 85.495 61.265 85.755 61.690 ;
        RECT 85.995 60.250 86.225 61.485 ;
        RECT 86.785 60.250 87.015 61.485 ;
        RECT 87.375 60.250 87.605 61.485 ;
        RECT 77.975 58.880 78.235 59.670 ;
        RECT 74.835 58.650 76.075 58.880 ;
        RECT 76.995 58.650 78.235 58.880 ;
        RECT 80.160 58.880 80.420 59.760 ;
        RECT 80.660 59.040 80.890 59.930 ;
        RECT 81.450 59.040 81.680 59.930 ;
        RECT 82.040 59.040 82.270 59.930 ;
        RECT 82.830 59.040 83.060 60.005 ;
        RECT 85.980 59.930 86.240 60.250 ;
        RECT 86.770 59.930 87.030 60.250 ;
        RECT 87.360 59.930 87.620 60.250 ;
        RECT 88.165 60.175 88.395 61.485 ;
        RECT 88.585 60.615 88.845 61.690 ;
        RECT 89.005 60.175 89.175 62.115 ;
        RECT 88.165 60.005 89.175 60.175 ;
        RECT 89.320 60.005 89.675 62.115 ;
        RECT 90.045 62.390 90.400 64.585 ;
        RECT 91.320 64.520 91.550 65.485 ;
        RECT 92.110 64.610 92.340 65.485 ;
        RECT 92.700 64.610 92.930 65.485 ;
        RECT 93.490 64.610 93.720 65.485 ;
        RECT 93.960 64.855 94.220 65.645 ;
        RECT 96.155 65.645 97.395 65.875 ;
        RECT 98.315 65.645 99.555 65.875 ;
        RECT 96.155 64.950 96.415 65.645 ;
        RECT 90.540 64.350 91.550 64.520 ;
        RECT 90.540 62.390 90.710 64.350 ;
        RECT 90.870 62.835 91.130 63.970 ;
        RECT 91.320 63.040 91.550 64.350 ;
        RECT 92.095 64.290 92.355 64.610 ;
        RECT 92.685 64.290 92.945 64.610 ;
        RECT 93.475 64.290 93.735 64.610 ;
        RECT 92.110 63.040 92.340 64.290 ;
        RECT 92.700 63.040 92.930 64.290 ;
        RECT 93.490 63.040 93.720 64.290 ;
        RECT 93.960 62.835 94.220 63.340 ;
        RECT 90.870 62.605 92.060 62.835 ;
        RECT 92.980 62.605 94.220 62.835 ;
        RECT 94.645 62.390 95.000 64.580 ;
        RECT 90.045 62.115 90.710 62.390 ;
        RECT 94.330 62.115 95.000 62.390 ;
        RECT 90.045 60.010 90.400 62.115 ;
        RECT 90.820 61.690 92.060 61.920 ;
        RECT 92.980 61.690 94.170 61.920 ;
        RECT 90.820 61.265 91.080 61.690 ;
        RECT 91.320 60.250 91.550 61.485 ;
        RECT 92.110 60.250 92.340 61.485 ;
        RECT 92.700 60.250 92.930 61.485 ;
        RECT 83.300 58.880 83.560 59.670 ;
        RECT 80.160 58.650 81.400 58.880 ;
        RECT 82.320 58.650 83.560 58.880 ;
        RECT 85.495 58.880 85.755 59.760 ;
        RECT 85.995 59.040 86.225 59.930 ;
        RECT 86.785 59.040 87.015 59.930 ;
        RECT 87.375 59.040 87.605 59.930 ;
        RECT 88.165 59.040 88.395 60.005 ;
        RECT 91.305 59.930 91.565 60.250 ;
        RECT 92.095 59.930 92.355 60.250 ;
        RECT 92.685 59.930 92.945 60.250 ;
        RECT 93.490 60.175 93.720 61.485 ;
        RECT 93.910 60.615 94.170 61.690 ;
        RECT 94.330 60.175 94.500 62.115 ;
        RECT 93.490 60.005 94.500 60.175 ;
        RECT 94.645 60.005 95.000 62.115 ;
        RECT 95.380 62.390 95.735 64.585 ;
        RECT 96.655 64.520 96.885 65.485 ;
        RECT 97.445 64.610 97.675 65.485 ;
        RECT 98.035 64.610 98.265 65.485 ;
        RECT 98.825 64.610 99.055 65.485 ;
        RECT 99.295 64.855 99.555 65.645 ;
        RECT 101.480 65.645 102.720 65.875 ;
        RECT 103.640 65.645 104.880 65.875 ;
        RECT 101.480 64.950 101.740 65.645 ;
        RECT 95.875 64.350 96.885 64.520 ;
        RECT 95.875 62.390 96.045 64.350 ;
        RECT 96.205 62.835 96.465 63.970 ;
        RECT 96.655 63.040 96.885 64.350 ;
        RECT 97.430 64.290 97.690 64.610 ;
        RECT 98.020 64.290 98.280 64.610 ;
        RECT 98.810 64.290 99.070 64.610 ;
        RECT 97.445 63.040 97.675 64.290 ;
        RECT 98.035 63.040 98.265 64.290 ;
        RECT 98.825 63.040 99.055 64.290 ;
        RECT 99.295 62.835 99.555 63.340 ;
        RECT 96.205 62.605 97.395 62.835 ;
        RECT 98.315 62.605 99.555 62.835 ;
        RECT 99.980 62.390 100.335 64.580 ;
        RECT 95.380 62.115 96.045 62.390 ;
        RECT 99.665 62.115 100.335 62.390 ;
        RECT 95.380 60.010 95.735 62.115 ;
        RECT 96.155 61.690 97.395 61.920 ;
        RECT 98.315 61.690 99.505 61.920 ;
        RECT 96.155 61.265 96.415 61.690 ;
        RECT 96.655 60.250 96.885 61.485 ;
        RECT 97.445 60.250 97.675 61.485 ;
        RECT 98.035 60.250 98.265 61.485 ;
        RECT 88.635 58.880 88.895 59.670 ;
        RECT 85.495 58.650 86.735 58.880 ;
        RECT 87.655 58.650 88.895 58.880 ;
        RECT 90.820 58.880 91.080 59.760 ;
        RECT 91.320 59.040 91.550 59.930 ;
        RECT 92.110 59.040 92.340 59.930 ;
        RECT 92.700 59.040 92.930 59.930 ;
        RECT 93.490 59.040 93.720 60.005 ;
        RECT 96.640 59.930 96.900 60.250 ;
        RECT 97.430 59.930 97.690 60.250 ;
        RECT 98.020 59.930 98.280 60.250 ;
        RECT 98.825 60.175 99.055 61.485 ;
        RECT 99.245 60.615 99.505 61.690 ;
        RECT 99.665 60.175 99.835 62.115 ;
        RECT 98.825 60.005 99.835 60.175 ;
        RECT 99.980 60.005 100.335 62.115 ;
        RECT 100.705 62.390 101.060 64.585 ;
        RECT 101.980 64.520 102.210 65.485 ;
        RECT 102.770 64.610 103.000 65.485 ;
        RECT 103.360 64.610 103.590 65.485 ;
        RECT 104.150 64.610 104.380 65.485 ;
        RECT 104.620 64.855 104.880 65.645 ;
        RECT 106.815 65.645 108.055 65.875 ;
        RECT 108.975 65.645 110.215 65.875 ;
        RECT 106.815 64.950 107.075 65.645 ;
        RECT 101.200 64.350 102.210 64.520 ;
        RECT 101.200 62.390 101.370 64.350 ;
        RECT 101.530 62.835 101.790 63.970 ;
        RECT 101.980 63.040 102.210 64.350 ;
        RECT 102.755 64.290 103.015 64.610 ;
        RECT 103.345 64.290 103.605 64.610 ;
        RECT 104.135 64.290 104.395 64.610 ;
        RECT 102.770 63.040 103.000 64.290 ;
        RECT 103.360 63.040 103.590 64.290 ;
        RECT 104.150 63.040 104.380 64.290 ;
        RECT 104.620 62.835 104.880 63.340 ;
        RECT 101.530 62.605 102.720 62.835 ;
        RECT 103.640 62.605 104.880 62.835 ;
        RECT 105.305 62.390 105.660 64.580 ;
        RECT 100.705 62.115 101.370 62.390 ;
        RECT 104.990 62.115 105.660 62.390 ;
        RECT 100.705 60.010 101.060 62.115 ;
        RECT 101.480 61.690 102.720 61.920 ;
        RECT 103.640 61.690 104.830 61.920 ;
        RECT 101.480 61.265 101.740 61.690 ;
        RECT 101.980 60.250 102.210 61.485 ;
        RECT 102.770 60.250 103.000 61.485 ;
        RECT 103.360 60.250 103.590 61.485 ;
        RECT 93.960 58.880 94.220 59.670 ;
        RECT 90.820 58.650 92.060 58.880 ;
        RECT 92.980 58.650 94.220 58.880 ;
        RECT 96.155 58.880 96.415 59.760 ;
        RECT 96.655 59.040 96.885 59.930 ;
        RECT 97.445 59.040 97.675 59.930 ;
        RECT 98.035 59.040 98.265 59.930 ;
        RECT 98.825 59.040 99.055 60.005 ;
        RECT 101.965 59.930 102.225 60.250 ;
        RECT 102.755 59.930 103.015 60.250 ;
        RECT 103.345 59.930 103.605 60.250 ;
        RECT 104.150 60.175 104.380 61.485 ;
        RECT 104.570 60.615 104.830 61.690 ;
        RECT 104.990 60.175 105.160 62.115 ;
        RECT 104.150 60.005 105.160 60.175 ;
        RECT 105.305 60.005 105.660 62.115 ;
        RECT 106.040 62.390 106.395 64.585 ;
        RECT 107.315 64.520 107.545 65.485 ;
        RECT 108.105 64.610 108.335 65.485 ;
        RECT 108.695 64.610 108.925 65.485 ;
        RECT 109.485 64.610 109.715 65.485 ;
        RECT 109.955 64.855 110.215 65.645 ;
        RECT 112.140 65.645 113.380 65.875 ;
        RECT 114.300 65.645 115.540 65.875 ;
        RECT 112.140 64.950 112.400 65.645 ;
        RECT 106.535 64.350 107.545 64.520 ;
        RECT 106.535 62.390 106.705 64.350 ;
        RECT 106.865 62.835 107.125 63.970 ;
        RECT 107.315 63.040 107.545 64.350 ;
        RECT 108.090 64.290 108.350 64.610 ;
        RECT 108.680 64.290 108.940 64.610 ;
        RECT 109.470 64.290 109.730 64.610 ;
        RECT 108.105 63.040 108.335 64.290 ;
        RECT 108.695 63.040 108.925 64.290 ;
        RECT 109.485 63.040 109.715 64.290 ;
        RECT 109.955 62.835 110.215 63.340 ;
        RECT 106.865 62.605 108.055 62.835 ;
        RECT 108.975 62.605 110.215 62.835 ;
        RECT 110.640 62.390 110.995 64.580 ;
        RECT 106.040 62.115 106.705 62.390 ;
        RECT 110.325 62.115 110.995 62.390 ;
        RECT 106.040 60.010 106.395 62.115 ;
        RECT 106.815 61.690 108.055 61.920 ;
        RECT 108.975 61.690 110.165 61.920 ;
        RECT 106.815 61.265 107.075 61.690 ;
        RECT 107.315 60.250 107.545 61.485 ;
        RECT 108.105 60.250 108.335 61.485 ;
        RECT 108.695 60.250 108.925 61.485 ;
        RECT 99.295 58.880 99.555 59.670 ;
        RECT 96.155 58.650 97.395 58.880 ;
        RECT 98.315 58.650 99.555 58.880 ;
        RECT 101.480 58.880 101.740 59.760 ;
        RECT 101.980 59.040 102.210 59.930 ;
        RECT 102.770 59.040 103.000 59.930 ;
        RECT 103.360 59.040 103.590 59.930 ;
        RECT 104.150 59.040 104.380 60.005 ;
        RECT 107.300 59.930 107.560 60.250 ;
        RECT 108.090 59.930 108.350 60.250 ;
        RECT 108.680 59.930 108.940 60.250 ;
        RECT 109.485 60.175 109.715 61.485 ;
        RECT 109.905 60.615 110.165 61.690 ;
        RECT 110.325 60.175 110.495 62.115 ;
        RECT 109.485 60.005 110.495 60.175 ;
        RECT 110.640 60.005 110.995 62.115 ;
        RECT 111.365 62.390 111.720 64.585 ;
        RECT 112.640 64.520 112.870 65.485 ;
        RECT 113.430 64.610 113.660 65.485 ;
        RECT 114.020 64.610 114.250 65.485 ;
        RECT 114.810 64.610 115.040 65.485 ;
        RECT 115.280 64.855 115.540 65.645 ;
        RECT 117.475 65.645 118.715 65.875 ;
        RECT 119.635 65.645 120.875 65.875 ;
        RECT 117.475 64.950 117.735 65.645 ;
        RECT 111.860 64.350 112.870 64.520 ;
        RECT 111.860 62.390 112.030 64.350 ;
        RECT 112.190 62.835 112.450 63.970 ;
        RECT 112.640 63.040 112.870 64.350 ;
        RECT 113.415 64.290 113.675 64.610 ;
        RECT 114.005 64.290 114.265 64.610 ;
        RECT 114.795 64.290 115.055 64.610 ;
        RECT 113.430 63.040 113.660 64.290 ;
        RECT 114.020 63.040 114.250 64.290 ;
        RECT 114.810 63.040 115.040 64.290 ;
        RECT 115.280 62.835 115.540 63.340 ;
        RECT 112.190 62.605 113.380 62.835 ;
        RECT 114.300 62.605 115.540 62.835 ;
        RECT 115.965 62.390 116.320 64.580 ;
        RECT 111.365 62.115 112.030 62.390 ;
        RECT 115.650 62.115 116.320 62.390 ;
        RECT 111.365 60.010 111.720 62.115 ;
        RECT 112.140 61.690 113.380 61.920 ;
        RECT 114.300 61.690 115.490 61.920 ;
        RECT 112.140 61.265 112.400 61.690 ;
        RECT 112.640 60.250 112.870 61.485 ;
        RECT 113.430 60.250 113.660 61.485 ;
        RECT 114.020 60.250 114.250 61.485 ;
        RECT 104.620 58.880 104.880 59.670 ;
        RECT 101.480 58.650 102.720 58.880 ;
        RECT 103.640 58.650 104.880 58.880 ;
        RECT 106.815 58.880 107.075 59.760 ;
        RECT 107.315 59.040 107.545 59.930 ;
        RECT 108.105 59.040 108.335 59.930 ;
        RECT 108.695 59.040 108.925 59.930 ;
        RECT 109.485 59.040 109.715 60.005 ;
        RECT 112.625 59.930 112.885 60.250 ;
        RECT 113.415 59.930 113.675 60.250 ;
        RECT 114.005 59.930 114.265 60.250 ;
        RECT 114.810 60.175 115.040 61.485 ;
        RECT 115.230 60.615 115.490 61.690 ;
        RECT 115.650 60.175 115.820 62.115 ;
        RECT 114.810 60.005 115.820 60.175 ;
        RECT 115.965 60.005 116.320 62.115 ;
        RECT 116.700 62.390 117.055 64.585 ;
        RECT 117.975 64.520 118.205 65.485 ;
        RECT 118.765 64.610 118.995 65.485 ;
        RECT 119.355 64.610 119.585 65.485 ;
        RECT 120.145 64.610 120.375 65.485 ;
        RECT 120.615 64.855 120.875 65.645 ;
        RECT 117.195 64.350 118.205 64.520 ;
        RECT 117.195 62.390 117.365 64.350 ;
        RECT 117.525 62.835 117.785 63.970 ;
        RECT 117.975 63.040 118.205 64.350 ;
        RECT 118.750 64.290 119.010 64.610 ;
        RECT 119.340 64.290 119.600 64.610 ;
        RECT 120.130 64.290 120.390 64.610 ;
        RECT 118.765 63.040 118.995 64.290 ;
        RECT 119.355 63.040 119.585 64.290 ;
        RECT 120.145 63.040 120.375 64.290 ;
        RECT 120.615 62.835 120.875 63.340 ;
        RECT 117.525 62.605 118.715 62.835 ;
        RECT 119.635 62.605 120.875 62.835 ;
        RECT 121.300 62.390 121.655 64.580 ;
        RECT 116.700 62.115 117.365 62.390 ;
        RECT 120.985 62.115 121.655 62.390 ;
        RECT 116.700 60.010 117.055 62.115 ;
        RECT 117.475 61.690 118.715 61.920 ;
        RECT 119.635 61.690 120.825 61.920 ;
        RECT 117.475 61.265 117.735 61.690 ;
        RECT 117.975 60.250 118.205 61.485 ;
        RECT 118.765 60.250 118.995 61.485 ;
        RECT 119.355 60.250 119.585 61.485 ;
        RECT 109.955 58.880 110.215 59.670 ;
        RECT 106.815 58.650 108.055 58.880 ;
        RECT 108.975 58.650 110.215 58.880 ;
        RECT 112.140 58.880 112.400 59.760 ;
        RECT 112.640 59.040 112.870 59.930 ;
        RECT 113.430 59.040 113.660 59.930 ;
        RECT 114.020 59.040 114.250 59.930 ;
        RECT 114.810 59.040 115.040 60.005 ;
        RECT 117.960 59.930 118.220 60.250 ;
        RECT 118.750 59.930 119.010 60.250 ;
        RECT 119.340 59.930 119.600 60.250 ;
        RECT 120.145 60.175 120.375 61.485 ;
        RECT 120.565 60.615 120.825 61.690 ;
        RECT 120.985 60.175 121.155 62.115 ;
        RECT 120.145 60.005 121.155 60.175 ;
        RECT 121.300 60.005 121.655 62.115 ;
        RECT 122.025 62.390 122.380 64.600 ;
        RECT 123.300 64.520 123.530 65.485 ;
        RECT 124.090 64.610 124.320 65.485 ;
        RECT 124.680 64.610 124.910 65.485 ;
        RECT 125.470 64.610 125.700 65.485 ;
        RECT 122.520 64.350 123.530 64.520 ;
        RECT 122.520 62.390 122.690 64.350 ;
        RECT 123.300 63.040 123.530 64.350 ;
        RECT 124.075 64.290 124.335 64.610 ;
        RECT 124.665 64.290 124.925 64.610 ;
        RECT 125.455 64.290 125.715 64.610 ;
        RECT 124.090 63.040 124.320 64.290 ;
        RECT 124.680 63.040 124.910 64.290 ;
        RECT 125.470 63.040 125.700 64.290 ;
        RECT 126.625 62.390 126.980 64.600 ;
        RECT 122.025 62.115 122.690 62.390 ;
        RECT 126.310 62.115 126.980 62.390 ;
        RECT 122.025 60.025 122.380 62.115 ;
        RECT 123.300 60.250 123.530 61.485 ;
        RECT 124.090 60.250 124.320 61.485 ;
        RECT 124.680 60.250 124.910 61.485 ;
        RECT 115.280 58.880 115.540 59.670 ;
        RECT 112.140 58.650 113.380 58.880 ;
        RECT 114.300 58.650 115.540 58.880 ;
        RECT 117.475 58.880 117.735 59.760 ;
        RECT 117.975 59.040 118.205 59.930 ;
        RECT 118.765 59.040 118.995 59.930 ;
        RECT 119.355 59.040 119.585 59.930 ;
        RECT 120.145 59.040 120.375 60.005 ;
        RECT 123.285 59.930 123.545 60.250 ;
        RECT 124.075 59.930 124.335 60.250 ;
        RECT 124.665 59.930 124.925 60.250 ;
        RECT 125.470 60.175 125.700 61.485 ;
        RECT 126.310 60.175 126.480 62.115 ;
        RECT 125.470 60.005 126.480 60.175 ;
        RECT 126.625 60.025 126.980 62.115 ;
        RECT 120.615 58.880 120.875 59.670 ;
        RECT 123.300 59.040 123.530 59.930 ;
        RECT 124.090 59.040 124.320 59.930 ;
        RECT 124.680 59.040 124.910 59.930 ;
        RECT 125.470 59.040 125.700 60.005 ;
        RECT 117.475 58.650 118.715 58.880 ;
        RECT 119.635 58.650 120.875 58.880 ;
        RECT 37.520 58.110 38.760 58.340 ;
        RECT 39.680 58.110 40.920 58.340 ;
        RECT 23.485 57.535 23.745 57.540 ;
        RECT 10.510 56.015 10.810 57.465 ;
        RECT 15.985 57.300 23.805 57.535 ;
        RECT 11.745 56.915 13.345 57.205 ;
        RECT 14.165 56.915 20.945 57.150 ;
        RECT 16.040 56.730 17.645 56.760 ;
        RECT 21.425 56.730 23.805 57.300 ;
        RECT 15.985 56.495 23.805 56.730 ;
        RECT 16.040 56.470 17.645 56.495 ;
        RECT 31.420 54.855 31.775 57.065 ;
        RECT 32.695 56.985 32.925 57.950 ;
        RECT 33.485 57.075 33.715 57.950 ;
        RECT 34.075 57.075 34.305 57.950 ;
        RECT 34.865 57.075 35.095 57.950 ;
        RECT 37.520 57.415 37.780 58.110 ;
        RECT 31.915 56.815 32.925 56.985 ;
        RECT 31.915 54.855 32.085 56.815 ;
        RECT 32.695 55.505 32.925 56.815 ;
        RECT 33.470 56.755 33.730 57.075 ;
        RECT 34.060 56.755 34.320 57.075 ;
        RECT 34.850 56.755 35.110 57.075 ;
        RECT 33.485 55.505 33.715 56.755 ;
        RECT 34.075 55.505 34.305 56.755 ;
        RECT 34.865 55.505 35.095 56.755 ;
        RECT 36.020 54.855 36.375 57.065 ;
        RECT 31.420 54.580 32.085 54.855 ;
        RECT 35.705 54.580 36.375 54.855 ;
        RECT 10.500 52.470 10.820 52.955 ;
        RECT 16.115 52.580 24.175 52.815 ;
        RECT 10.500 52.140 11.960 52.470 ;
        RECT 10.500 51.920 10.820 52.140 ;
        RECT 12.400 51.395 12.720 52.385 ;
        RECT 14.585 52.140 16.005 52.465 ;
        RECT 19.990 52.010 24.175 52.580 ;
        RECT 31.420 52.490 31.775 54.580 ;
        RECT 32.695 52.715 32.925 53.950 ;
        RECT 33.485 52.715 33.715 53.950 ;
        RECT 34.075 52.715 34.305 53.950 ;
        RECT 32.680 52.395 32.940 52.715 ;
        RECT 33.470 52.395 33.730 52.715 ;
        RECT 34.060 52.395 34.320 52.715 ;
        RECT 34.865 52.640 35.095 53.950 ;
        RECT 35.705 52.640 35.875 54.580 ;
        RECT 34.865 52.470 35.875 52.640 ;
        RECT 36.020 52.490 36.375 54.580 ;
        RECT 36.745 54.855 37.100 57.050 ;
        RECT 38.020 56.985 38.250 57.950 ;
        RECT 38.810 57.075 39.040 57.950 ;
        RECT 39.400 57.075 39.630 57.950 ;
        RECT 40.190 57.075 40.420 57.950 ;
        RECT 40.660 57.320 40.920 58.110 ;
        RECT 42.855 58.110 44.095 58.340 ;
        RECT 45.015 58.110 46.255 58.340 ;
        RECT 42.855 57.415 43.115 58.110 ;
        RECT 37.240 56.815 38.250 56.985 ;
        RECT 37.240 54.855 37.410 56.815 ;
        RECT 37.570 55.300 37.830 56.435 ;
        RECT 38.020 55.505 38.250 56.815 ;
        RECT 38.795 56.755 39.055 57.075 ;
        RECT 39.385 56.755 39.645 57.075 ;
        RECT 40.175 56.755 40.435 57.075 ;
        RECT 38.810 55.505 39.040 56.755 ;
        RECT 39.400 55.505 39.630 56.755 ;
        RECT 40.190 55.505 40.420 56.755 ;
        RECT 40.660 55.300 40.920 55.805 ;
        RECT 37.570 55.070 38.760 55.300 ;
        RECT 39.680 55.070 40.920 55.300 ;
        RECT 41.345 54.855 41.700 57.045 ;
        RECT 36.745 54.580 37.410 54.855 ;
        RECT 41.030 54.580 41.700 54.855 ;
        RECT 36.745 52.475 37.100 54.580 ;
        RECT 37.520 54.155 38.760 54.385 ;
        RECT 39.680 54.155 40.870 54.385 ;
        RECT 37.520 53.730 37.780 54.155 ;
        RECT 38.020 52.715 38.250 53.950 ;
        RECT 38.810 52.715 39.040 53.950 ;
        RECT 39.400 52.715 39.630 53.950 ;
        RECT 16.115 51.775 24.175 52.010 ;
        RECT 32.695 51.505 32.925 52.395 ;
        RECT 33.485 51.505 33.715 52.395 ;
        RECT 34.075 51.505 34.305 52.395 ;
        RECT 34.865 51.505 35.095 52.470 ;
        RECT 38.005 52.395 38.265 52.715 ;
        RECT 38.795 52.395 39.055 52.715 ;
        RECT 39.385 52.395 39.645 52.715 ;
        RECT 40.190 52.640 40.420 53.950 ;
        RECT 40.610 53.080 40.870 54.155 ;
        RECT 41.030 52.640 41.200 54.580 ;
        RECT 40.190 52.470 41.200 52.640 ;
        RECT 41.345 52.470 41.700 54.580 ;
        RECT 42.080 54.855 42.435 57.050 ;
        RECT 43.355 56.985 43.585 57.950 ;
        RECT 44.145 57.075 44.375 57.950 ;
        RECT 44.735 57.075 44.965 57.950 ;
        RECT 45.525 57.075 45.755 57.950 ;
        RECT 45.995 57.320 46.255 58.110 ;
        RECT 48.180 58.110 49.420 58.340 ;
        RECT 50.340 58.110 51.580 58.340 ;
        RECT 48.180 57.415 48.440 58.110 ;
        RECT 42.575 56.815 43.585 56.985 ;
        RECT 42.575 54.855 42.745 56.815 ;
        RECT 42.905 55.300 43.165 56.435 ;
        RECT 43.355 55.505 43.585 56.815 ;
        RECT 44.130 56.755 44.390 57.075 ;
        RECT 44.720 56.755 44.980 57.075 ;
        RECT 45.510 56.755 45.770 57.075 ;
        RECT 44.145 55.505 44.375 56.755 ;
        RECT 44.735 55.505 44.965 56.755 ;
        RECT 45.525 55.505 45.755 56.755 ;
        RECT 45.995 55.300 46.255 55.805 ;
        RECT 42.905 55.070 44.095 55.300 ;
        RECT 45.015 55.070 46.255 55.300 ;
        RECT 46.680 54.855 47.035 57.045 ;
        RECT 42.080 54.580 42.745 54.855 ;
        RECT 46.365 54.580 47.035 54.855 ;
        RECT 42.080 52.475 42.435 54.580 ;
        RECT 42.855 54.155 44.095 54.385 ;
        RECT 45.015 54.155 46.205 54.385 ;
        RECT 42.855 53.730 43.115 54.155 ;
        RECT 43.355 52.715 43.585 53.950 ;
        RECT 44.145 52.715 44.375 53.950 ;
        RECT 44.735 52.715 44.965 53.950 ;
        RECT 12.425 51.380 12.715 51.395 ;
        RECT 37.520 51.345 37.780 52.225 ;
        RECT 38.020 51.505 38.250 52.395 ;
        RECT 38.810 51.505 39.040 52.395 ;
        RECT 39.400 51.505 39.630 52.395 ;
        RECT 40.190 51.505 40.420 52.470 ;
        RECT 43.340 52.395 43.600 52.715 ;
        RECT 44.130 52.395 44.390 52.715 ;
        RECT 44.720 52.395 44.980 52.715 ;
        RECT 45.525 52.640 45.755 53.950 ;
        RECT 45.945 53.080 46.205 54.155 ;
        RECT 46.365 52.640 46.535 54.580 ;
        RECT 45.525 52.470 46.535 52.640 ;
        RECT 46.680 52.470 47.035 54.580 ;
        RECT 47.405 54.855 47.760 57.050 ;
        RECT 48.680 56.985 48.910 57.950 ;
        RECT 49.470 57.075 49.700 57.950 ;
        RECT 50.060 57.075 50.290 57.950 ;
        RECT 50.850 57.075 51.080 57.950 ;
        RECT 51.320 57.320 51.580 58.110 ;
        RECT 53.515 58.110 54.755 58.340 ;
        RECT 55.675 58.110 56.915 58.340 ;
        RECT 53.515 57.415 53.775 58.110 ;
        RECT 47.900 56.815 48.910 56.985 ;
        RECT 47.900 54.855 48.070 56.815 ;
        RECT 48.230 55.300 48.490 56.435 ;
        RECT 48.680 55.505 48.910 56.815 ;
        RECT 49.455 56.755 49.715 57.075 ;
        RECT 50.045 56.755 50.305 57.075 ;
        RECT 50.835 56.755 51.095 57.075 ;
        RECT 49.470 55.505 49.700 56.755 ;
        RECT 50.060 55.505 50.290 56.755 ;
        RECT 50.850 55.505 51.080 56.755 ;
        RECT 51.320 55.300 51.580 55.805 ;
        RECT 48.230 55.070 49.420 55.300 ;
        RECT 50.340 55.070 51.580 55.300 ;
        RECT 52.005 54.855 52.360 57.045 ;
        RECT 47.405 54.580 48.070 54.855 ;
        RECT 51.690 54.580 52.360 54.855 ;
        RECT 47.405 52.475 47.760 54.580 ;
        RECT 48.180 54.155 49.420 54.385 ;
        RECT 50.340 54.155 51.530 54.385 ;
        RECT 48.180 53.730 48.440 54.155 ;
        RECT 48.680 52.715 48.910 53.950 ;
        RECT 49.470 52.715 49.700 53.950 ;
        RECT 50.060 52.715 50.290 53.950 ;
        RECT 40.660 51.345 40.920 52.135 ;
        RECT 37.520 51.115 38.760 51.345 ;
        RECT 39.680 51.115 40.920 51.345 ;
        RECT 42.855 51.345 43.115 52.225 ;
        RECT 43.355 51.505 43.585 52.395 ;
        RECT 44.145 51.505 44.375 52.395 ;
        RECT 44.735 51.505 44.965 52.395 ;
        RECT 45.525 51.505 45.755 52.470 ;
        RECT 48.665 52.395 48.925 52.715 ;
        RECT 49.455 52.395 49.715 52.715 ;
        RECT 50.045 52.395 50.305 52.715 ;
        RECT 50.850 52.640 51.080 53.950 ;
        RECT 51.270 53.080 51.530 54.155 ;
        RECT 51.690 52.640 51.860 54.580 ;
        RECT 50.850 52.470 51.860 52.640 ;
        RECT 52.005 52.470 52.360 54.580 ;
        RECT 52.740 54.855 53.095 57.050 ;
        RECT 54.015 56.985 54.245 57.950 ;
        RECT 54.805 57.075 55.035 57.950 ;
        RECT 55.395 57.075 55.625 57.950 ;
        RECT 56.185 57.075 56.415 57.950 ;
        RECT 56.655 57.320 56.915 58.110 ;
        RECT 58.840 58.110 60.080 58.340 ;
        RECT 61.000 58.110 62.240 58.340 ;
        RECT 58.840 57.415 59.100 58.110 ;
        RECT 53.235 56.815 54.245 56.985 ;
        RECT 53.235 54.855 53.405 56.815 ;
        RECT 53.565 55.300 53.825 56.435 ;
        RECT 54.015 55.505 54.245 56.815 ;
        RECT 54.790 56.755 55.050 57.075 ;
        RECT 55.380 56.755 55.640 57.075 ;
        RECT 56.170 56.755 56.430 57.075 ;
        RECT 54.805 55.505 55.035 56.755 ;
        RECT 55.395 55.505 55.625 56.755 ;
        RECT 56.185 55.505 56.415 56.755 ;
        RECT 56.655 55.300 56.915 55.805 ;
        RECT 53.565 55.070 54.755 55.300 ;
        RECT 55.675 55.070 56.915 55.300 ;
        RECT 57.340 54.855 57.695 57.045 ;
        RECT 52.740 54.580 53.405 54.855 ;
        RECT 57.025 54.580 57.695 54.855 ;
        RECT 52.740 52.475 53.095 54.580 ;
        RECT 53.515 54.155 54.755 54.385 ;
        RECT 55.675 54.155 56.865 54.385 ;
        RECT 53.515 53.730 53.775 54.155 ;
        RECT 54.015 52.715 54.245 53.950 ;
        RECT 54.805 52.715 55.035 53.950 ;
        RECT 55.395 52.715 55.625 53.950 ;
        RECT 45.995 51.345 46.255 52.135 ;
        RECT 42.855 51.115 44.095 51.345 ;
        RECT 45.015 51.115 46.255 51.345 ;
        RECT 48.180 51.345 48.440 52.225 ;
        RECT 48.680 51.505 48.910 52.395 ;
        RECT 49.470 51.505 49.700 52.395 ;
        RECT 50.060 51.505 50.290 52.395 ;
        RECT 50.850 51.505 51.080 52.470 ;
        RECT 54.000 52.395 54.260 52.715 ;
        RECT 54.790 52.395 55.050 52.715 ;
        RECT 55.380 52.395 55.640 52.715 ;
        RECT 56.185 52.640 56.415 53.950 ;
        RECT 56.605 53.080 56.865 54.155 ;
        RECT 57.025 52.640 57.195 54.580 ;
        RECT 56.185 52.470 57.195 52.640 ;
        RECT 57.340 52.470 57.695 54.580 ;
        RECT 58.065 54.855 58.420 57.050 ;
        RECT 59.340 56.985 59.570 57.950 ;
        RECT 60.130 57.075 60.360 57.950 ;
        RECT 60.720 57.075 60.950 57.950 ;
        RECT 61.510 57.075 61.740 57.950 ;
        RECT 61.980 57.320 62.240 58.110 ;
        RECT 64.175 58.110 65.415 58.340 ;
        RECT 66.335 58.110 67.575 58.340 ;
        RECT 64.175 57.415 64.435 58.110 ;
        RECT 58.560 56.815 59.570 56.985 ;
        RECT 58.560 54.855 58.730 56.815 ;
        RECT 58.890 55.300 59.150 56.435 ;
        RECT 59.340 55.505 59.570 56.815 ;
        RECT 60.115 56.755 60.375 57.075 ;
        RECT 60.705 56.755 60.965 57.075 ;
        RECT 61.495 56.755 61.755 57.075 ;
        RECT 60.130 55.505 60.360 56.755 ;
        RECT 60.720 55.505 60.950 56.755 ;
        RECT 61.510 55.505 61.740 56.755 ;
        RECT 61.980 55.300 62.240 55.805 ;
        RECT 58.890 55.070 60.080 55.300 ;
        RECT 61.000 55.070 62.240 55.300 ;
        RECT 62.665 54.855 63.020 57.045 ;
        RECT 58.065 54.580 58.730 54.855 ;
        RECT 62.350 54.580 63.020 54.855 ;
        RECT 58.065 52.475 58.420 54.580 ;
        RECT 58.840 54.155 60.080 54.385 ;
        RECT 61.000 54.155 62.190 54.385 ;
        RECT 58.840 53.730 59.100 54.155 ;
        RECT 59.340 52.715 59.570 53.950 ;
        RECT 60.130 52.715 60.360 53.950 ;
        RECT 60.720 52.715 60.950 53.950 ;
        RECT 51.320 51.345 51.580 52.135 ;
        RECT 48.180 51.115 49.420 51.345 ;
        RECT 50.340 51.115 51.580 51.345 ;
        RECT 53.515 51.345 53.775 52.225 ;
        RECT 54.015 51.505 54.245 52.395 ;
        RECT 54.805 51.505 55.035 52.395 ;
        RECT 55.395 51.505 55.625 52.395 ;
        RECT 56.185 51.505 56.415 52.470 ;
        RECT 59.325 52.395 59.585 52.715 ;
        RECT 60.115 52.395 60.375 52.715 ;
        RECT 60.705 52.395 60.965 52.715 ;
        RECT 61.510 52.640 61.740 53.950 ;
        RECT 61.930 53.080 62.190 54.155 ;
        RECT 62.350 52.640 62.520 54.580 ;
        RECT 61.510 52.470 62.520 52.640 ;
        RECT 62.665 52.470 63.020 54.580 ;
        RECT 63.400 54.855 63.755 57.050 ;
        RECT 64.675 56.985 64.905 57.950 ;
        RECT 65.465 57.075 65.695 57.950 ;
        RECT 66.055 57.075 66.285 57.950 ;
        RECT 66.845 57.075 67.075 57.950 ;
        RECT 67.315 57.320 67.575 58.110 ;
        RECT 69.500 58.110 70.740 58.340 ;
        RECT 71.660 58.110 72.900 58.340 ;
        RECT 69.500 57.415 69.760 58.110 ;
        RECT 63.895 56.815 64.905 56.985 ;
        RECT 63.895 54.855 64.065 56.815 ;
        RECT 64.225 55.300 64.485 56.435 ;
        RECT 64.675 55.505 64.905 56.815 ;
        RECT 65.450 56.755 65.710 57.075 ;
        RECT 66.040 56.755 66.300 57.075 ;
        RECT 66.830 56.755 67.090 57.075 ;
        RECT 65.465 55.505 65.695 56.755 ;
        RECT 66.055 55.505 66.285 56.755 ;
        RECT 66.845 55.505 67.075 56.755 ;
        RECT 67.315 55.300 67.575 55.805 ;
        RECT 64.225 55.070 65.415 55.300 ;
        RECT 66.335 55.070 67.575 55.300 ;
        RECT 68.000 54.855 68.355 57.045 ;
        RECT 63.400 54.580 64.065 54.855 ;
        RECT 67.685 54.580 68.355 54.855 ;
        RECT 63.400 52.475 63.755 54.580 ;
        RECT 64.175 54.155 65.415 54.385 ;
        RECT 66.335 54.155 67.525 54.385 ;
        RECT 64.175 53.730 64.435 54.155 ;
        RECT 64.675 52.715 64.905 53.950 ;
        RECT 65.465 52.715 65.695 53.950 ;
        RECT 66.055 52.715 66.285 53.950 ;
        RECT 56.655 51.345 56.915 52.135 ;
        RECT 53.515 51.115 54.755 51.345 ;
        RECT 55.675 51.115 56.915 51.345 ;
        RECT 58.840 51.345 59.100 52.225 ;
        RECT 59.340 51.505 59.570 52.395 ;
        RECT 60.130 51.505 60.360 52.395 ;
        RECT 60.720 51.505 60.950 52.395 ;
        RECT 61.510 51.505 61.740 52.470 ;
        RECT 64.660 52.395 64.920 52.715 ;
        RECT 65.450 52.395 65.710 52.715 ;
        RECT 66.040 52.395 66.300 52.715 ;
        RECT 66.845 52.640 67.075 53.950 ;
        RECT 67.265 53.080 67.525 54.155 ;
        RECT 67.685 52.640 67.855 54.580 ;
        RECT 66.845 52.470 67.855 52.640 ;
        RECT 68.000 52.470 68.355 54.580 ;
        RECT 68.725 54.855 69.080 57.050 ;
        RECT 70.000 56.985 70.230 57.950 ;
        RECT 70.790 57.075 71.020 57.950 ;
        RECT 71.380 57.075 71.610 57.950 ;
        RECT 72.170 57.075 72.400 57.950 ;
        RECT 72.640 57.320 72.900 58.110 ;
        RECT 74.835 58.110 76.075 58.340 ;
        RECT 76.995 58.110 78.235 58.340 ;
        RECT 74.835 57.415 75.095 58.110 ;
        RECT 69.220 56.815 70.230 56.985 ;
        RECT 69.220 54.855 69.390 56.815 ;
        RECT 69.550 55.300 69.810 56.435 ;
        RECT 70.000 55.505 70.230 56.815 ;
        RECT 70.775 56.755 71.035 57.075 ;
        RECT 71.365 56.755 71.625 57.075 ;
        RECT 72.155 56.755 72.415 57.075 ;
        RECT 70.790 55.505 71.020 56.755 ;
        RECT 71.380 55.505 71.610 56.755 ;
        RECT 72.170 55.505 72.400 56.755 ;
        RECT 72.640 55.300 72.900 55.805 ;
        RECT 69.550 55.070 70.740 55.300 ;
        RECT 71.660 55.070 72.900 55.300 ;
        RECT 73.325 54.855 73.680 57.045 ;
        RECT 68.725 54.580 69.390 54.855 ;
        RECT 73.010 54.580 73.680 54.855 ;
        RECT 68.725 52.475 69.080 54.580 ;
        RECT 69.500 54.155 70.740 54.385 ;
        RECT 71.660 54.155 72.850 54.385 ;
        RECT 69.500 53.730 69.760 54.155 ;
        RECT 70.000 52.715 70.230 53.950 ;
        RECT 70.790 52.715 71.020 53.950 ;
        RECT 71.380 52.715 71.610 53.950 ;
        RECT 61.980 51.345 62.240 52.135 ;
        RECT 58.840 51.115 60.080 51.345 ;
        RECT 61.000 51.115 62.240 51.345 ;
        RECT 64.175 51.345 64.435 52.225 ;
        RECT 64.675 51.505 64.905 52.395 ;
        RECT 65.465 51.505 65.695 52.395 ;
        RECT 66.055 51.505 66.285 52.395 ;
        RECT 66.845 51.505 67.075 52.470 ;
        RECT 69.985 52.395 70.245 52.715 ;
        RECT 70.775 52.395 71.035 52.715 ;
        RECT 71.365 52.395 71.625 52.715 ;
        RECT 72.170 52.640 72.400 53.950 ;
        RECT 72.590 53.080 72.850 54.155 ;
        RECT 73.010 52.640 73.180 54.580 ;
        RECT 72.170 52.470 73.180 52.640 ;
        RECT 73.325 52.470 73.680 54.580 ;
        RECT 74.060 54.855 74.415 57.050 ;
        RECT 75.335 56.985 75.565 57.950 ;
        RECT 76.125 57.075 76.355 57.950 ;
        RECT 76.715 57.075 76.945 57.950 ;
        RECT 77.505 57.075 77.735 57.950 ;
        RECT 77.975 57.320 78.235 58.110 ;
        RECT 80.160 58.110 81.400 58.340 ;
        RECT 82.320 58.110 83.560 58.340 ;
        RECT 80.160 57.415 80.420 58.110 ;
        RECT 74.555 56.815 75.565 56.985 ;
        RECT 74.555 54.855 74.725 56.815 ;
        RECT 74.885 55.300 75.145 56.435 ;
        RECT 75.335 55.505 75.565 56.815 ;
        RECT 76.110 56.755 76.370 57.075 ;
        RECT 76.700 56.755 76.960 57.075 ;
        RECT 77.490 56.755 77.750 57.075 ;
        RECT 76.125 55.505 76.355 56.755 ;
        RECT 76.715 55.505 76.945 56.755 ;
        RECT 77.505 55.505 77.735 56.755 ;
        RECT 77.975 55.300 78.235 55.805 ;
        RECT 74.885 55.070 76.075 55.300 ;
        RECT 76.995 55.070 78.235 55.300 ;
        RECT 78.660 54.855 79.015 57.045 ;
        RECT 74.060 54.580 74.725 54.855 ;
        RECT 78.345 54.580 79.015 54.855 ;
        RECT 74.060 52.475 74.415 54.580 ;
        RECT 74.835 54.155 76.075 54.385 ;
        RECT 76.995 54.155 78.185 54.385 ;
        RECT 74.835 53.730 75.095 54.155 ;
        RECT 75.335 52.715 75.565 53.950 ;
        RECT 76.125 52.715 76.355 53.950 ;
        RECT 76.715 52.715 76.945 53.950 ;
        RECT 67.315 51.345 67.575 52.135 ;
        RECT 64.175 51.115 65.415 51.345 ;
        RECT 66.335 51.115 67.575 51.345 ;
        RECT 69.500 51.345 69.760 52.225 ;
        RECT 70.000 51.505 70.230 52.395 ;
        RECT 70.790 51.505 71.020 52.395 ;
        RECT 71.380 51.505 71.610 52.395 ;
        RECT 72.170 51.505 72.400 52.470 ;
        RECT 75.320 52.395 75.580 52.715 ;
        RECT 76.110 52.395 76.370 52.715 ;
        RECT 76.700 52.395 76.960 52.715 ;
        RECT 77.505 52.640 77.735 53.950 ;
        RECT 77.925 53.080 78.185 54.155 ;
        RECT 78.345 52.640 78.515 54.580 ;
        RECT 77.505 52.470 78.515 52.640 ;
        RECT 78.660 52.470 79.015 54.580 ;
        RECT 79.385 54.855 79.740 57.050 ;
        RECT 80.660 56.985 80.890 57.950 ;
        RECT 81.450 57.075 81.680 57.950 ;
        RECT 82.040 57.075 82.270 57.950 ;
        RECT 82.830 57.075 83.060 57.950 ;
        RECT 83.300 57.320 83.560 58.110 ;
        RECT 85.495 58.110 86.735 58.340 ;
        RECT 87.655 58.110 88.895 58.340 ;
        RECT 85.495 57.415 85.755 58.110 ;
        RECT 79.880 56.815 80.890 56.985 ;
        RECT 79.880 54.855 80.050 56.815 ;
        RECT 80.210 55.300 80.470 56.435 ;
        RECT 80.660 55.505 80.890 56.815 ;
        RECT 81.435 56.755 81.695 57.075 ;
        RECT 82.025 56.755 82.285 57.075 ;
        RECT 82.815 56.755 83.075 57.075 ;
        RECT 81.450 55.505 81.680 56.755 ;
        RECT 82.040 55.505 82.270 56.755 ;
        RECT 82.830 55.505 83.060 56.755 ;
        RECT 83.300 55.300 83.560 55.805 ;
        RECT 80.210 55.070 81.400 55.300 ;
        RECT 82.320 55.070 83.560 55.300 ;
        RECT 83.985 54.855 84.340 57.045 ;
        RECT 79.385 54.580 80.050 54.855 ;
        RECT 83.670 54.580 84.340 54.855 ;
        RECT 79.385 52.475 79.740 54.580 ;
        RECT 80.160 54.155 81.400 54.385 ;
        RECT 82.320 54.155 83.510 54.385 ;
        RECT 80.160 53.730 80.420 54.155 ;
        RECT 80.660 52.715 80.890 53.950 ;
        RECT 81.450 52.715 81.680 53.950 ;
        RECT 82.040 52.715 82.270 53.950 ;
        RECT 72.640 51.345 72.900 52.135 ;
        RECT 69.500 51.115 70.740 51.345 ;
        RECT 71.660 51.115 72.900 51.345 ;
        RECT 74.835 51.345 75.095 52.225 ;
        RECT 75.335 51.505 75.565 52.395 ;
        RECT 76.125 51.505 76.355 52.395 ;
        RECT 76.715 51.505 76.945 52.395 ;
        RECT 77.505 51.505 77.735 52.470 ;
        RECT 80.645 52.395 80.905 52.715 ;
        RECT 81.435 52.395 81.695 52.715 ;
        RECT 82.025 52.395 82.285 52.715 ;
        RECT 82.830 52.640 83.060 53.950 ;
        RECT 83.250 53.080 83.510 54.155 ;
        RECT 83.670 52.640 83.840 54.580 ;
        RECT 82.830 52.470 83.840 52.640 ;
        RECT 83.985 52.470 84.340 54.580 ;
        RECT 84.720 54.855 85.075 57.050 ;
        RECT 85.995 56.985 86.225 57.950 ;
        RECT 86.785 57.075 87.015 57.950 ;
        RECT 87.375 57.075 87.605 57.950 ;
        RECT 88.165 57.075 88.395 57.950 ;
        RECT 88.635 57.320 88.895 58.110 ;
        RECT 90.820 58.110 92.060 58.340 ;
        RECT 92.980 58.110 94.220 58.340 ;
        RECT 90.820 57.415 91.080 58.110 ;
        RECT 85.215 56.815 86.225 56.985 ;
        RECT 85.215 54.855 85.385 56.815 ;
        RECT 85.545 55.300 85.805 56.435 ;
        RECT 85.995 55.505 86.225 56.815 ;
        RECT 86.770 56.755 87.030 57.075 ;
        RECT 87.360 56.755 87.620 57.075 ;
        RECT 88.150 56.755 88.410 57.075 ;
        RECT 86.785 55.505 87.015 56.755 ;
        RECT 87.375 55.505 87.605 56.755 ;
        RECT 88.165 55.505 88.395 56.755 ;
        RECT 88.635 55.300 88.895 55.805 ;
        RECT 85.545 55.070 86.735 55.300 ;
        RECT 87.655 55.070 88.895 55.300 ;
        RECT 89.320 54.855 89.675 57.045 ;
        RECT 84.720 54.580 85.385 54.855 ;
        RECT 89.005 54.580 89.675 54.855 ;
        RECT 84.720 52.475 85.075 54.580 ;
        RECT 85.495 54.155 86.735 54.385 ;
        RECT 87.655 54.155 88.845 54.385 ;
        RECT 85.495 53.730 85.755 54.155 ;
        RECT 85.995 52.715 86.225 53.950 ;
        RECT 86.785 52.715 87.015 53.950 ;
        RECT 87.375 52.715 87.605 53.950 ;
        RECT 77.975 51.345 78.235 52.135 ;
        RECT 74.835 51.115 76.075 51.345 ;
        RECT 76.995 51.115 78.235 51.345 ;
        RECT 80.160 51.345 80.420 52.225 ;
        RECT 80.660 51.505 80.890 52.395 ;
        RECT 81.450 51.505 81.680 52.395 ;
        RECT 82.040 51.505 82.270 52.395 ;
        RECT 82.830 51.505 83.060 52.470 ;
        RECT 85.980 52.395 86.240 52.715 ;
        RECT 86.770 52.395 87.030 52.715 ;
        RECT 87.360 52.395 87.620 52.715 ;
        RECT 88.165 52.640 88.395 53.950 ;
        RECT 88.585 53.080 88.845 54.155 ;
        RECT 89.005 52.640 89.175 54.580 ;
        RECT 88.165 52.470 89.175 52.640 ;
        RECT 89.320 52.470 89.675 54.580 ;
        RECT 90.045 54.855 90.400 57.050 ;
        RECT 91.320 56.985 91.550 57.950 ;
        RECT 92.110 57.075 92.340 57.950 ;
        RECT 92.700 57.075 92.930 57.950 ;
        RECT 93.490 57.075 93.720 57.950 ;
        RECT 93.960 57.320 94.220 58.110 ;
        RECT 96.155 58.110 97.395 58.340 ;
        RECT 98.315 58.110 99.555 58.340 ;
        RECT 96.155 57.415 96.415 58.110 ;
        RECT 90.540 56.815 91.550 56.985 ;
        RECT 90.540 54.855 90.710 56.815 ;
        RECT 90.870 55.300 91.130 56.435 ;
        RECT 91.320 55.505 91.550 56.815 ;
        RECT 92.095 56.755 92.355 57.075 ;
        RECT 92.685 56.755 92.945 57.075 ;
        RECT 93.475 56.755 93.735 57.075 ;
        RECT 92.110 55.505 92.340 56.755 ;
        RECT 92.700 55.505 92.930 56.755 ;
        RECT 93.490 55.505 93.720 56.755 ;
        RECT 93.960 55.300 94.220 55.805 ;
        RECT 90.870 55.070 92.060 55.300 ;
        RECT 92.980 55.070 94.220 55.300 ;
        RECT 94.645 54.855 95.000 57.045 ;
        RECT 90.045 54.580 90.710 54.855 ;
        RECT 94.330 54.580 95.000 54.855 ;
        RECT 90.045 52.475 90.400 54.580 ;
        RECT 90.820 54.155 92.060 54.385 ;
        RECT 92.980 54.155 94.170 54.385 ;
        RECT 90.820 53.730 91.080 54.155 ;
        RECT 91.320 52.715 91.550 53.950 ;
        RECT 92.110 52.715 92.340 53.950 ;
        RECT 92.700 52.715 92.930 53.950 ;
        RECT 83.300 51.345 83.560 52.135 ;
        RECT 80.160 51.115 81.400 51.345 ;
        RECT 82.320 51.115 83.560 51.345 ;
        RECT 85.495 51.345 85.755 52.225 ;
        RECT 85.995 51.505 86.225 52.395 ;
        RECT 86.785 51.505 87.015 52.395 ;
        RECT 87.375 51.505 87.605 52.395 ;
        RECT 88.165 51.505 88.395 52.470 ;
        RECT 91.305 52.395 91.565 52.715 ;
        RECT 92.095 52.395 92.355 52.715 ;
        RECT 92.685 52.395 92.945 52.715 ;
        RECT 93.490 52.640 93.720 53.950 ;
        RECT 93.910 53.080 94.170 54.155 ;
        RECT 94.330 52.640 94.500 54.580 ;
        RECT 93.490 52.470 94.500 52.640 ;
        RECT 94.645 52.470 95.000 54.580 ;
        RECT 95.380 54.855 95.735 57.050 ;
        RECT 96.655 56.985 96.885 57.950 ;
        RECT 97.445 57.075 97.675 57.950 ;
        RECT 98.035 57.075 98.265 57.950 ;
        RECT 98.825 57.075 99.055 57.950 ;
        RECT 99.295 57.320 99.555 58.110 ;
        RECT 101.480 58.110 102.720 58.340 ;
        RECT 103.640 58.110 104.880 58.340 ;
        RECT 101.480 57.415 101.740 58.110 ;
        RECT 95.875 56.815 96.885 56.985 ;
        RECT 95.875 54.855 96.045 56.815 ;
        RECT 96.205 55.300 96.465 56.435 ;
        RECT 96.655 55.505 96.885 56.815 ;
        RECT 97.430 56.755 97.690 57.075 ;
        RECT 98.020 56.755 98.280 57.075 ;
        RECT 98.810 56.755 99.070 57.075 ;
        RECT 97.445 55.505 97.675 56.755 ;
        RECT 98.035 55.505 98.265 56.755 ;
        RECT 98.825 55.505 99.055 56.755 ;
        RECT 99.295 55.300 99.555 55.805 ;
        RECT 96.205 55.070 97.395 55.300 ;
        RECT 98.315 55.070 99.555 55.300 ;
        RECT 99.980 54.855 100.335 57.045 ;
        RECT 95.380 54.580 96.045 54.855 ;
        RECT 99.665 54.580 100.335 54.855 ;
        RECT 95.380 52.475 95.735 54.580 ;
        RECT 96.155 54.155 97.395 54.385 ;
        RECT 98.315 54.155 99.505 54.385 ;
        RECT 96.155 53.730 96.415 54.155 ;
        RECT 96.655 52.715 96.885 53.950 ;
        RECT 97.445 52.715 97.675 53.950 ;
        RECT 98.035 52.715 98.265 53.950 ;
        RECT 88.635 51.345 88.895 52.135 ;
        RECT 85.495 51.115 86.735 51.345 ;
        RECT 87.655 51.115 88.895 51.345 ;
        RECT 90.820 51.345 91.080 52.225 ;
        RECT 91.320 51.505 91.550 52.395 ;
        RECT 92.110 51.505 92.340 52.395 ;
        RECT 92.700 51.505 92.930 52.395 ;
        RECT 93.490 51.505 93.720 52.470 ;
        RECT 96.640 52.395 96.900 52.715 ;
        RECT 97.430 52.395 97.690 52.715 ;
        RECT 98.020 52.395 98.280 52.715 ;
        RECT 98.825 52.640 99.055 53.950 ;
        RECT 99.245 53.080 99.505 54.155 ;
        RECT 99.665 52.640 99.835 54.580 ;
        RECT 98.825 52.470 99.835 52.640 ;
        RECT 99.980 52.470 100.335 54.580 ;
        RECT 100.705 54.855 101.060 57.050 ;
        RECT 101.980 56.985 102.210 57.950 ;
        RECT 102.770 57.075 103.000 57.950 ;
        RECT 103.360 57.075 103.590 57.950 ;
        RECT 104.150 57.075 104.380 57.950 ;
        RECT 104.620 57.320 104.880 58.110 ;
        RECT 106.815 58.110 108.055 58.340 ;
        RECT 108.975 58.110 110.215 58.340 ;
        RECT 106.815 57.415 107.075 58.110 ;
        RECT 101.200 56.815 102.210 56.985 ;
        RECT 101.200 54.855 101.370 56.815 ;
        RECT 101.530 55.300 101.790 56.435 ;
        RECT 101.980 55.505 102.210 56.815 ;
        RECT 102.755 56.755 103.015 57.075 ;
        RECT 103.345 56.755 103.605 57.075 ;
        RECT 104.135 56.755 104.395 57.075 ;
        RECT 102.770 55.505 103.000 56.755 ;
        RECT 103.360 55.505 103.590 56.755 ;
        RECT 104.150 55.505 104.380 56.755 ;
        RECT 104.620 55.300 104.880 55.805 ;
        RECT 101.530 55.070 102.720 55.300 ;
        RECT 103.640 55.070 104.880 55.300 ;
        RECT 105.305 54.855 105.660 57.045 ;
        RECT 100.705 54.580 101.370 54.855 ;
        RECT 104.990 54.580 105.660 54.855 ;
        RECT 100.705 52.475 101.060 54.580 ;
        RECT 101.480 54.155 102.720 54.385 ;
        RECT 103.640 54.155 104.830 54.385 ;
        RECT 101.480 53.730 101.740 54.155 ;
        RECT 101.980 52.715 102.210 53.950 ;
        RECT 102.770 52.715 103.000 53.950 ;
        RECT 103.360 52.715 103.590 53.950 ;
        RECT 93.960 51.345 94.220 52.135 ;
        RECT 90.820 51.115 92.060 51.345 ;
        RECT 92.980 51.115 94.220 51.345 ;
        RECT 96.155 51.345 96.415 52.225 ;
        RECT 96.655 51.505 96.885 52.395 ;
        RECT 97.445 51.505 97.675 52.395 ;
        RECT 98.035 51.505 98.265 52.395 ;
        RECT 98.825 51.505 99.055 52.470 ;
        RECT 101.965 52.395 102.225 52.715 ;
        RECT 102.755 52.395 103.015 52.715 ;
        RECT 103.345 52.395 103.605 52.715 ;
        RECT 104.150 52.640 104.380 53.950 ;
        RECT 104.570 53.080 104.830 54.155 ;
        RECT 104.990 52.640 105.160 54.580 ;
        RECT 104.150 52.470 105.160 52.640 ;
        RECT 105.305 52.470 105.660 54.580 ;
        RECT 106.040 54.855 106.395 57.050 ;
        RECT 107.315 56.985 107.545 57.950 ;
        RECT 108.105 57.075 108.335 57.950 ;
        RECT 108.695 57.075 108.925 57.950 ;
        RECT 109.485 57.075 109.715 57.950 ;
        RECT 109.955 57.320 110.215 58.110 ;
        RECT 112.140 58.110 113.380 58.340 ;
        RECT 114.300 58.110 115.540 58.340 ;
        RECT 112.140 57.415 112.400 58.110 ;
        RECT 106.535 56.815 107.545 56.985 ;
        RECT 106.535 54.855 106.705 56.815 ;
        RECT 106.865 55.300 107.125 56.435 ;
        RECT 107.315 55.505 107.545 56.815 ;
        RECT 108.090 56.755 108.350 57.075 ;
        RECT 108.680 56.755 108.940 57.075 ;
        RECT 109.470 56.755 109.730 57.075 ;
        RECT 108.105 55.505 108.335 56.755 ;
        RECT 108.695 55.505 108.925 56.755 ;
        RECT 109.485 55.505 109.715 56.755 ;
        RECT 109.955 55.300 110.215 55.805 ;
        RECT 106.865 55.070 108.055 55.300 ;
        RECT 108.975 55.070 110.215 55.300 ;
        RECT 110.640 54.855 110.995 57.045 ;
        RECT 106.040 54.580 106.705 54.855 ;
        RECT 110.325 54.580 110.995 54.855 ;
        RECT 106.040 52.475 106.395 54.580 ;
        RECT 106.815 54.155 108.055 54.385 ;
        RECT 108.975 54.155 110.165 54.385 ;
        RECT 106.815 53.730 107.075 54.155 ;
        RECT 107.315 52.715 107.545 53.950 ;
        RECT 108.105 52.715 108.335 53.950 ;
        RECT 108.695 52.715 108.925 53.950 ;
        RECT 99.295 51.345 99.555 52.135 ;
        RECT 96.155 51.115 97.395 51.345 ;
        RECT 98.315 51.115 99.555 51.345 ;
        RECT 101.480 51.345 101.740 52.225 ;
        RECT 101.980 51.505 102.210 52.395 ;
        RECT 102.770 51.505 103.000 52.395 ;
        RECT 103.360 51.505 103.590 52.395 ;
        RECT 104.150 51.505 104.380 52.470 ;
        RECT 107.300 52.395 107.560 52.715 ;
        RECT 108.090 52.395 108.350 52.715 ;
        RECT 108.680 52.395 108.940 52.715 ;
        RECT 109.485 52.640 109.715 53.950 ;
        RECT 109.905 53.080 110.165 54.155 ;
        RECT 110.325 52.640 110.495 54.580 ;
        RECT 109.485 52.470 110.495 52.640 ;
        RECT 110.640 52.470 110.995 54.580 ;
        RECT 111.365 54.855 111.720 57.050 ;
        RECT 112.640 56.985 112.870 57.950 ;
        RECT 113.430 57.075 113.660 57.950 ;
        RECT 114.020 57.075 114.250 57.950 ;
        RECT 114.810 57.075 115.040 57.950 ;
        RECT 115.280 57.320 115.540 58.110 ;
        RECT 117.475 58.110 118.715 58.340 ;
        RECT 119.635 58.110 120.875 58.340 ;
        RECT 117.475 57.415 117.735 58.110 ;
        RECT 111.860 56.815 112.870 56.985 ;
        RECT 111.860 54.855 112.030 56.815 ;
        RECT 112.190 55.300 112.450 56.435 ;
        RECT 112.640 55.505 112.870 56.815 ;
        RECT 113.415 56.755 113.675 57.075 ;
        RECT 114.005 56.755 114.265 57.075 ;
        RECT 114.795 56.755 115.055 57.075 ;
        RECT 113.430 55.505 113.660 56.755 ;
        RECT 114.020 55.505 114.250 56.755 ;
        RECT 114.810 55.505 115.040 56.755 ;
        RECT 115.280 55.300 115.540 55.805 ;
        RECT 112.190 55.070 113.380 55.300 ;
        RECT 114.300 55.070 115.540 55.300 ;
        RECT 115.965 54.855 116.320 57.045 ;
        RECT 111.365 54.580 112.030 54.855 ;
        RECT 115.650 54.580 116.320 54.855 ;
        RECT 111.365 52.475 111.720 54.580 ;
        RECT 112.140 54.155 113.380 54.385 ;
        RECT 114.300 54.155 115.490 54.385 ;
        RECT 112.140 53.730 112.400 54.155 ;
        RECT 112.640 52.715 112.870 53.950 ;
        RECT 113.430 52.715 113.660 53.950 ;
        RECT 114.020 52.715 114.250 53.950 ;
        RECT 104.620 51.345 104.880 52.135 ;
        RECT 101.480 51.115 102.720 51.345 ;
        RECT 103.640 51.115 104.880 51.345 ;
        RECT 106.815 51.345 107.075 52.225 ;
        RECT 107.315 51.505 107.545 52.395 ;
        RECT 108.105 51.505 108.335 52.395 ;
        RECT 108.695 51.505 108.925 52.395 ;
        RECT 109.485 51.505 109.715 52.470 ;
        RECT 112.625 52.395 112.885 52.715 ;
        RECT 113.415 52.395 113.675 52.715 ;
        RECT 114.005 52.395 114.265 52.715 ;
        RECT 114.810 52.640 115.040 53.950 ;
        RECT 115.230 53.080 115.490 54.155 ;
        RECT 115.650 52.640 115.820 54.580 ;
        RECT 114.810 52.470 115.820 52.640 ;
        RECT 115.965 52.470 116.320 54.580 ;
        RECT 116.700 54.855 117.055 57.050 ;
        RECT 117.975 56.985 118.205 57.950 ;
        RECT 118.765 57.075 118.995 57.950 ;
        RECT 119.355 57.075 119.585 57.950 ;
        RECT 120.145 57.075 120.375 57.950 ;
        RECT 120.615 57.320 120.875 58.110 ;
        RECT 117.195 56.815 118.205 56.985 ;
        RECT 117.195 54.855 117.365 56.815 ;
        RECT 117.525 55.300 117.785 56.435 ;
        RECT 117.975 55.505 118.205 56.815 ;
        RECT 118.750 56.755 119.010 57.075 ;
        RECT 119.340 56.755 119.600 57.075 ;
        RECT 120.130 56.755 120.390 57.075 ;
        RECT 118.765 55.505 118.995 56.755 ;
        RECT 119.355 55.505 119.585 56.755 ;
        RECT 120.145 55.505 120.375 56.755 ;
        RECT 120.615 55.300 120.875 55.805 ;
        RECT 117.525 55.070 118.715 55.300 ;
        RECT 119.635 55.070 120.875 55.300 ;
        RECT 121.300 54.855 121.655 57.045 ;
        RECT 116.700 54.580 117.365 54.855 ;
        RECT 120.985 54.580 121.655 54.855 ;
        RECT 116.700 52.475 117.055 54.580 ;
        RECT 117.475 54.155 118.715 54.385 ;
        RECT 119.635 54.155 120.825 54.385 ;
        RECT 117.475 53.730 117.735 54.155 ;
        RECT 117.975 52.715 118.205 53.950 ;
        RECT 118.765 52.715 118.995 53.950 ;
        RECT 119.355 52.715 119.585 53.950 ;
        RECT 109.955 51.345 110.215 52.135 ;
        RECT 106.815 51.115 108.055 51.345 ;
        RECT 108.975 51.115 110.215 51.345 ;
        RECT 112.140 51.345 112.400 52.225 ;
        RECT 112.640 51.505 112.870 52.395 ;
        RECT 113.430 51.505 113.660 52.395 ;
        RECT 114.020 51.505 114.250 52.395 ;
        RECT 114.810 51.505 115.040 52.470 ;
        RECT 117.960 52.395 118.220 52.715 ;
        RECT 118.750 52.395 119.010 52.715 ;
        RECT 119.340 52.395 119.600 52.715 ;
        RECT 120.145 52.640 120.375 53.950 ;
        RECT 120.565 53.080 120.825 54.155 ;
        RECT 120.985 52.640 121.155 54.580 ;
        RECT 120.145 52.470 121.155 52.640 ;
        RECT 121.300 52.470 121.655 54.580 ;
        RECT 122.025 54.855 122.380 57.065 ;
        RECT 123.300 56.985 123.530 57.950 ;
        RECT 124.090 57.075 124.320 57.950 ;
        RECT 124.680 57.075 124.910 57.950 ;
        RECT 125.470 57.075 125.700 57.950 ;
        RECT 122.520 56.815 123.530 56.985 ;
        RECT 122.520 54.855 122.690 56.815 ;
        RECT 123.300 55.505 123.530 56.815 ;
        RECT 124.075 56.755 124.335 57.075 ;
        RECT 124.665 56.755 124.925 57.075 ;
        RECT 125.455 56.755 125.715 57.075 ;
        RECT 124.090 55.505 124.320 56.755 ;
        RECT 124.680 55.505 124.910 56.755 ;
        RECT 125.470 55.505 125.700 56.755 ;
        RECT 126.625 54.855 126.980 57.065 ;
        RECT 122.025 54.580 122.690 54.855 ;
        RECT 126.310 54.580 126.980 54.855 ;
        RECT 122.025 52.490 122.380 54.580 ;
        RECT 123.300 52.715 123.530 53.950 ;
        RECT 124.090 52.715 124.320 53.950 ;
        RECT 124.680 52.715 124.910 53.950 ;
        RECT 115.280 51.345 115.540 52.135 ;
        RECT 112.140 51.115 113.380 51.345 ;
        RECT 114.300 51.115 115.540 51.345 ;
        RECT 117.475 51.345 117.735 52.225 ;
        RECT 117.975 51.505 118.205 52.395 ;
        RECT 118.765 51.505 118.995 52.395 ;
        RECT 119.355 51.505 119.585 52.395 ;
        RECT 120.145 51.505 120.375 52.470 ;
        RECT 123.285 52.395 123.545 52.715 ;
        RECT 124.075 52.395 124.335 52.715 ;
        RECT 124.665 52.395 124.925 52.715 ;
        RECT 125.470 52.640 125.700 53.950 ;
        RECT 126.310 52.640 126.480 54.580 ;
        RECT 125.470 52.470 126.480 52.640 ;
        RECT 126.625 52.490 126.980 54.580 ;
        RECT 120.615 51.345 120.875 52.135 ;
        RECT 123.300 51.505 123.530 52.395 ;
        RECT 124.090 51.505 124.320 52.395 ;
        RECT 124.680 51.505 124.910 52.395 ;
        RECT 125.470 51.505 125.700 52.470 ;
        RECT 117.475 51.115 118.715 51.345 ;
        RECT 119.635 51.115 120.875 51.345 ;
        RECT 37.520 50.575 38.760 50.805 ;
        RECT 39.680 50.575 40.920 50.805 ;
        RECT 24.625 49.395 24.885 49.400 ;
        RECT 10.510 47.875 10.810 49.325 ;
        RECT 15.985 49.160 24.930 49.395 ;
        RECT 11.745 48.775 13.345 49.065 ;
        RECT 14.165 48.775 20.945 49.010 ;
        RECT 16.040 48.590 17.645 48.620 ;
        RECT 21.425 48.590 24.930 49.160 ;
        RECT 15.985 48.355 24.930 48.590 ;
        RECT 16.040 48.330 17.645 48.355 ;
        RECT 31.420 47.320 31.775 49.530 ;
        RECT 32.695 49.450 32.925 50.415 ;
        RECT 33.485 49.540 33.715 50.415 ;
        RECT 34.075 49.540 34.305 50.415 ;
        RECT 34.865 49.540 35.095 50.415 ;
        RECT 37.520 49.880 37.780 50.575 ;
        RECT 31.915 49.280 32.925 49.450 ;
        RECT 31.915 47.320 32.085 49.280 ;
        RECT 32.695 47.970 32.925 49.280 ;
        RECT 33.470 49.220 33.730 49.540 ;
        RECT 34.060 49.220 34.320 49.540 ;
        RECT 34.850 49.220 35.110 49.540 ;
        RECT 33.485 47.970 33.715 49.220 ;
        RECT 34.075 47.970 34.305 49.220 ;
        RECT 34.865 47.970 35.095 49.220 ;
        RECT 36.020 47.320 36.375 49.530 ;
        RECT 31.420 47.045 32.085 47.320 ;
        RECT 35.705 47.045 36.375 47.320 ;
        RECT 31.420 44.955 31.775 47.045 ;
        RECT 32.695 45.180 32.925 46.415 ;
        RECT 33.485 45.180 33.715 46.415 ;
        RECT 34.075 45.180 34.305 46.415 ;
        RECT 32.680 44.860 32.940 45.180 ;
        RECT 33.470 44.860 33.730 45.180 ;
        RECT 34.060 44.860 34.320 45.180 ;
        RECT 34.865 45.105 35.095 46.415 ;
        RECT 35.705 45.105 35.875 47.045 ;
        RECT 34.865 44.935 35.875 45.105 ;
        RECT 36.020 44.955 36.375 47.045 ;
        RECT 36.745 47.320 37.100 49.515 ;
        RECT 38.020 49.450 38.250 50.415 ;
        RECT 38.810 49.540 39.040 50.415 ;
        RECT 39.400 49.540 39.630 50.415 ;
        RECT 40.190 49.540 40.420 50.415 ;
        RECT 40.660 49.785 40.920 50.575 ;
        RECT 42.855 50.575 44.095 50.805 ;
        RECT 45.015 50.575 46.255 50.805 ;
        RECT 42.855 49.880 43.115 50.575 ;
        RECT 37.240 49.280 38.250 49.450 ;
        RECT 37.240 47.320 37.410 49.280 ;
        RECT 37.570 47.765 37.830 48.900 ;
        RECT 38.020 47.970 38.250 49.280 ;
        RECT 38.795 49.220 39.055 49.540 ;
        RECT 39.385 49.220 39.645 49.540 ;
        RECT 40.175 49.220 40.435 49.540 ;
        RECT 38.810 47.970 39.040 49.220 ;
        RECT 39.400 47.970 39.630 49.220 ;
        RECT 40.190 47.970 40.420 49.220 ;
        RECT 40.660 47.765 40.920 48.270 ;
        RECT 37.570 47.535 38.760 47.765 ;
        RECT 39.680 47.535 40.920 47.765 ;
        RECT 41.345 47.320 41.700 49.510 ;
        RECT 36.745 47.045 37.410 47.320 ;
        RECT 41.030 47.045 41.700 47.320 ;
        RECT 36.745 44.940 37.100 47.045 ;
        RECT 37.520 46.620 38.760 46.850 ;
        RECT 39.680 46.620 40.870 46.850 ;
        RECT 37.520 46.195 37.780 46.620 ;
        RECT 38.020 45.180 38.250 46.415 ;
        RECT 38.810 45.180 39.040 46.415 ;
        RECT 39.400 45.180 39.630 46.415 ;
        RECT 10.500 44.330 10.820 44.815 ;
        RECT 16.115 44.440 24.565 44.675 ;
        RECT 10.500 44.000 11.960 44.330 ;
        RECT 10.500 43.780 10.820 44.000 ;
        RECT 12.400 43.255 12.720 44.245 ;
        RECT 14.585 44.000 16.005 44.325 ;
        RECT 19.990 43.870 24.565 44.440 ;
        RECT 32.695 43.970 32.925 44.860 ;
        RECT 33.485 43.970 33.715 44.860 ;
        RECT 34.075 43.970 34.305 44.860 ;
        RECT 34.865 43.970 35.095 44.935 ;
        RECT 38.005 44.860 38.265 45.180 ;
        RECT 38.795 44.860 39.055 45.180 ;
        RECT 39.385 44.860 39.645 45.180 ;
        RECT 40.190 45.105 40.420 46.415 ;
        RECT 40.610 45.545 40.870 46.620 ;
        RECT 41.030 45.105 41.200 47.045 ;
        RECT 40.190 44.935 41.200 45.105 ;
        RECT 41.345 44.935 41.700 47.045 ;
        RECT 42.080 47.320 42.435 49.515 ;
        RECT 43.355 49.450 43.585 50.415 ;
        RECT 44.145 49.540 44.375 50.415 ;
        RECT 44.735 49.540 44.965 50.415 ;
        RECT 45.525 49.540 45.755 50.415 ;
        RECT 45.995 49.785 46.255 50.575 ;
        RECT 48.180 50.575 49.420 50.805 ;
        RECT 50.340 50.575 51.580 50.805 ;
        RECT 48.180 49.880 48.440 50.575 ;
        RECT 42.575 49.280 43.585 49.450 ;
        RECT 42.575 47.320 42.745 49.280 ;
        RECT 42.905 47.765 43.165 48.900 ;
        RECT 43.355 47.970 43.585 49.280 ;
        RECT 44.130 49.220 44.390 49.540 ;
        RECT 44.720 49.220 44.980 49.540 ;
        RECT 45.510 49.220 45.770 49.540 ;
        RECT 44.145 47.970 44.375 49.220 ;
        RECT 44.735 47.970 44.965 49.220 ;
        RECT 45.525 47.970 45.755 49.220 ;
        RECT 45.995 47.765 46.255 48.270 ;
        RECT 42.905 47.535 44.095 47.765 ;
        RECT 45.015 47.535 46.255 47.765 ;
        RECT 46.680 47.320 47.035 49.510 ;
        RECT 42.080 47.045 42.745 47.320 ;
        RECT 46.365 47.045 47.035 47.320 ;
        RECT 42.080 44.940 42.435 47.045 ;
        RECT 42.855 46.620 44.095 46.850 ;
        RECT 45.015 46.620 46.205 46.850 ;
        RECT 42.855 46.195 43.115 46.620 ;
        RECT 43.355 45.180 43.585 46.415 ;
        RECT 44.145 45.180 44.375 46.415 ;
        RECT 44.735 45.180 44.965 46.415 ;
        RECT 16.115 43.635 24.565 43.870 ;
        RECT 37.520 43.810 37.780 44.690 ;
        RECT 38.020 43.970 38.250 44.860 ;
        RECT 38.810 43.970 39.040 44.860 ;
        RECT 39.400 43.970 39.630 44.860 ;
        RECT 40.190 43.970 40.420 44.935 ;
        RECT 43.340 44.860 43.600 45.180 ;
        RECT 44.130 44.860 44.390 45.180 ;
        RECT 44.720 44.860 44.980 45.180 ;
        RECT 45.525 45.105 45.755 46.415 ;
        RECT 45.945 45.545 46.205 46.620 ;
        RECT 46.365 45.105 46.535 47.045 ;
        RECT 45.525 44.935 46.535 45.105 ;
        RECT 46.680 44.935 47.035 47.045 ;
        RECT 47.405 47.320 47.760 49.515 ;
        RECT 48.680 49.450 48.910 50.415 ;
        RECT 49.470 49.540 49.700 50.415 ;
        RECT 50.060 49.540 50.290 50.415 ;
        RECT 50.850 49.540 51.080 50.415 ;
        RECT 51.320 49.785 51.580 50.575 ;
        RECT 53.515 50.575 54.755 50.805 ;
        RECT 55.675 50.575 56.915 50.805 ;
        RECT 53.515 49.880 53.775 50.575 ;
        RECT 47.900 49.280 48.910 49.450 ;
        RECT 47.900 47.320 48.070 49.280 ;
        RECT 48.230 47.765 48.490 48.900 ;
        RECT 48.680 47.970 48.910 49.280 ;
        RECT 49.455 49.220 49.715 49.540 ;
        RECT 50.045 49.220 50.305 49.540 ;
        RECT 50.835 49.220 51.095 49.540 ;
        RECT 49.470 47.970 49.700 49.220 ;
        RECT 50.060 47.970 50.290 49.220 ;
        RECT 50.850 47.970 51.080 49.220 ;
        RECT 51.320 47.765 51.580 48.270 ;
        RECT 48.230 47.535 49.420 47.765 ;
        RECT 50.340 47.535 51.580 47.765 ;
        RECT 52.005 47.320 52.360 49.510 ;
        RECT 47.405 47.045 48.070 47.320 ;
        RECT 51.690 47.045 52.360 47.320 ;
        RECT 47.405 44.940 47.760 47.045 ;
        RECT 48.180 46.620 49.420 46.850 ;
        RECT 50.340 46.620 51.530 46.850 ;
        RECT 48.180 46.195 48.440 46.620 ;
        RECT 48.680 45.180 48.910 46.415 ;
        RECT 49.470 45.180 49.700 46.415 ;
        RECT 50.060 45.180 50.290 46.415 ;
        RECT 40.660 43.810 40.920 44.600 ;
        RECT 37.520 43.580 38.760 43.810 ;
        RECT 39.680 43.580 40.920 43.810 ;
        RECT 42.855 43.810 43.115 44.690 ;
        RECT 43.355 43.970 43.585 44.860 ;
        RECT 44.145 43.970 44.375 44.860 ;
        RECT 44.735 43.970 44.965 44.860 ;
        RECT 45.525 43.970 45.755 44.935 ;
        RECT 48.665 44.860 48.925 45.180 ;
        RECT 49.455 44.860 49.715 45.180 ;
        RECT 50.045 44.860 50.305 45.180 ;
        RECT 50.850 45.105 51.080 46.415 ;
        RECT 51.270 45.545 51.530 46.620 ;
        RECT 51.690 45.105 51.860 47.045 ;
        RECT 50.850 44.935 51.860 45.105 ;
        RECT 52.005 44.935 52.360 47.045 ;
        RECT 52.740 47.320 53.095 49.515 ;
        RECT 54.015 49.450 54.245 50.415 ;
        RECT 54.805 49.540 55.035 50.415 ;
        RECT 55.395 49.540 55.625 50.415 ;
        RECT 56.185 49.540 56.415 50.415 ;
        RECT 56.655 49.785 56.915 50.575 ;
        RECT 58.840 50.575 60.080 50.805 ;
        RECT 61.000 50.575 62.240 50.805 ;
        RECT 58.840 49.880 59.100 50.575 ;
        RECT 53.235 49.280 54.245 49.450 ;
        RECT 53.235 47.320 53.405 49.280 ;
        RECT 53.565 47.765 53.825 48.900 ;
        RECT 54.015 47.970 54.245 49.280 ;
        RECT 54.790 49.220 55.050 49.540 ;
        RECT 55.380 49.220 55.640 49.540 ;
        RECT 56.170 49.220 56.430 49.540 ;
        RECT 54.805 47.970 55.035 49.220 ;
        RECT 55.395 47.970 55.625 49.220 ;
        RECT 56.185 47.970 56.415 49.220 ;
        RECT 56.655 47.765 56.915 48.270 ;
        RECT 53.565 47.535 54.755 47.765 ;
        RECT 55.675 47.535 56.915 47.765 ;
        RECT 57.340 47.320 57.695 49.510 ;
        RECT 52.740 47.045 53.405 47.320 ;
        RECT 57.025 47.045 57.695 47.320 ;
        RECT 52.740 44.940 53.095 47.045 ;
        RECT 53.515 46.620 54.755 46.850 ;
        RECT 55.675 46.620 56.865 46.850 ;
        RECT 53.515 46.195 53.775 46.620 ;
        RECT 54.015 45.180 54.245 46.415 ;
        RECT 54.805 45.180 55.035 46.415 ;
        RECT 55.395 45.180 55.625 46.415 ;
        RECT 45.995 43.810 46.255 44.600 ;
        RECT 42.855 43.580 44.095 43.810 ;
        RECT 45.015 43.580 46.255 43.810 ;
        RECT 48.180 43.810 48.440 44.690 ;
        RECT 48.680 43.970 48.910 44.860 ;
        RECT 49.470 43.970 49.700 44.860 ;
        RECT 50.060 43.970 50.290 44.860 ;
        RECT 50.850 43.970 51.080 44.935 ;
        RECT 54.000 44.860 54.260 45.180 ;
        RECT 54.790 44.860 55.050 45.180 ;
        RECT 55.380 44.860 55.640 45.180 ;
        RECT 56.185 45.105 56.415 46.415 ;
        RECT 56.605 45.545 56.865 46.620 ;
        RECT 57.025 45.105 57.195 47.045 ;
        RECT 56.185 44.935 57.195 45.105 ;
        RECT 57.340 44.935 57.695 47.045 ;
        RECT 58.065 47.320 58.420 49.515 ;
        RECT 59.340 49.450 59.570 50.415 ;
        RECT 60.130 49.540 60.360 50.415 ;
        RECT 60.720 49.540 60.950 50.415 ;
        RECT 61.510 49.540 61.740 50.415 ;
        RECT 61.980 49.785 62.240 50.575 ;
        RECT 64.175 50.575 65.415 50.805 ;
        RECT 66.335 50.575 67.575 50.805 ;
        RECT 64.175 49.880 64.435 50.575 ;
        RECT 58.560 49.280 59.570 49.450 ;
        RECT 58.560 47.320 58.730 49.280 ;
        RECT 58.890 47.765 59.150 48.900 ;
        RECT 59.340 47.970 59.570 49.280 ;
        RECT 60.115 49.220 60.375 49.540 ;
        RECT 60.705 49.220 60.965 49.540 ;
        RECT 61.495 49.220 61.755 49.540 ;
        RECT 60.130 47.970 60.360 49.220 ;
        RECT 60.720 47.970 60.950 49.220 ;
        RECT 61.510 47.970 61.740 49.220 ;
        RECT 61.980 47.765 62.240 48.270 ;
        RECT 58.890 47.535 60.080 47.765 ;
        RECT 61.000 47.535 62.240 47.765 ;
        RECT 62.665 47.320 63.020 49.510 ;
        RECT 58.065 47.045 58.730 47.320 ;
        RECT 62.350 47.045 63.020 47.320 ;
        RECT 58.065 44.940 58.420 47.045 ;
        RECT 58.840 46.620 60.080 46.850 ;
        RECT 61.000 46.620 62.190 46.850 ;
        RECT 58.840 46.195 59.100 46.620 ;
        RECT 59.340 45.180 59.570 46.415 ;
        RECT 60.130 45.180 60.360 46.415 ;
        RECT 60.720 45.180 60.950 46.415 ;
        RECT 51.320 43.810 51.580 44.600 ;
        RECT 48.180 43.580 49.420 43.810 ;
        RECT 50.340 43.580 51.580 43.810 ;
        RECT 53.515 43.810 53.775 44.690 ;
        RECT 54.015 43.970 54.245 44.860 ;
        RECT 54.805 43.970 55.035 44.860 ;
        RECT 55.395 43.970 55.625 44.860 ;
        RECT 56.185 43.970 56.415 44.935 ;
        RECT 59.325 44.860 59.585 45.180 ;
        RECT 60.115 44.860 60.375 45.180 ;
        RECT 60.705 44.860 60.965 45.180 ;
        RECT 61.510 45.105 61.740 46.415 ;
        RECT 61.930 45.545 62.190 46.620 ;
        RECT 62.350 45.105 62.520 47.045 ;
        RECT 61.510 44.935 62.520 45.105 ;
        RECT 62.665 44.935 63.020 47.045 ;
        RECT 63.400 47.320 63.755 49.515 ;
        RECT 64.675 49.450 64.905 50.415 ;
        RECT 65.465 49.540 65.695 50.415 ;
        RECT 66.055 49.540 66.285 50.415 ;
        RECT 66.845 49.540 67.075 50.415 ;
        RECT 67.315 49.785 67.575 50.575 ;
        RECT 69.500 50.575 70.740 50.805 ;
        RECT 71.660 50.575 72.900 50.805 ;
        RECT 69.500 49.880 69.760 50.575 ;
        RECT 63.895 49.280 64.905 49.450 ;
        RECT 63.895 47.320 64.065 49.280 ;
        RECT 64.225 47.765 64.485 48.900 ;
        RECT 64.675 47.970 64.905 49.280 ;
        RECT 65.450 49.220 65.710 49.540 ;
        RECT 66.040 49.220 66.300 49.540 ;
        RECT 66.830 49.220 67.090 49.540 ;
        RECT 65.465 47.970 65.695 49.220 ;
        RECT 66.055 47.970 66.285 49.220 ;
        RECT 66.845 47.970 67.075 49.220 ;
        RECT 67.315 47.765 67.575 48.270 ;
        RECT 64.225 47.535 65.415 47.765 ;
        RECT 66.335 47.535 67.575 47.765 ;
        RECT 68.000 47.320 68.355 49.510 ;
        RECT 63.400 47.045 64.065 47.320 ;
        RECT 67.685 47.045 68.355 47.320 ;
        RECT 63.400 44.940 63.755 47.045 ;
        RECT 64.175 46.620 65.415 46.850 ;
        RECT 66.335 46.620 67.525 46.850 ;
        RECT 64.175 46.195 64.435 46.620 ;
        RECT 64.675 45.180 64.905 46.415 ;
        RECT 65.465 45.180 65.695 46.415 ;
        RECT 66.055 45.180 66.285 46.415 ;
        RECT 56.655 43.810 56.915 44.600 ;
        RECT 53.515 43.580 54.755 43.810 ;
        RECT 55.675 43.580 56.915 43.810 ;
        RECT 58.840 43.810 59.100 44.690 ;
        RECT 59.340 43.970 59.570 44.860 ;
        RECT 60.130 43.970 60.360 44.860 ;
        RECT 60.720 43.970 60.950 44.860 ;
        RECT 61.510 43.970 61.740 44.935 ;
        RECT 64.660 44.860 64.920 45.180 ;
        RECT 65.450 44.860 65.710 45.180 ;
        RECT 66.040 44.860 66.300 45.180 ;
        RECT 66.845 45.105 67.075 46.415 ;
        RECT 67.265 45.545 67.525 46.620 ;
        RECT 67.685 45.105 67.855 47.045 ;
        RECT 66.845 44.935 67.855 45.105 ;
        RECT 68.000 44.935 68.355 47.045 ;
        RECT 68.725 47.320 69.080 49.515 ;
        RECT 70.000 49.450 70.230 50.415 ;
        RECT 70.790 49.540 71.020 50.415 ;
        RECT 71.380 49.540 71.610 50.415 ;
        RECT 72.170 49.540 72.400 50.415 ;
        RECT 72.640 49.785 72.900 50.575 ;
        RECT 74.835 50.575 76.075 50.805 ;
        RECT 76.995 50.575 78.235 50.805 ;
        RECT 74.835 49.880 75.095 50.575 ;
        RECT 69.220 49.280 70.230 49.450 ;
        RECT 69.220 47.320 69.390 49.280 ;
        RECT 69.550 47.765 69.810 48.900 ;
        RECT 70.000 47.970 70.230 49.280 ;
        RECT 70.775 49.220 71.035 49.540 ;
        RECT 71.365 49.220 71.625 49.540 ;
        RECT 72.155 49.220 72.415 49.540 ;
        RECT 70.790 47.970 71.020 49.220 ;
        RECT 71.380 47.970 71.610 49.220 ;
        RECT 72.170 47.970 72.400 49.220 ;
        RECT 72.640 47.765 72.900 48.270 ;
        RECT 69.550 47.535 70.740 47.765 ;
        RECT 71.660 47.535 72.900 47.765 ;
        RECT 73.325 47.320 73.680 49.510 ;
        RECT 68.725 47.045 69.390 47.320 ;
        RECT 73.010 47.045 73.680 47.320 ;
        RECT 68.725 44.940 69.080 47.045 ;
        RECT 69.500 46.620 70.740 46.850 ;
        RECT 71.660 46.620 72.850 46.850 ;
        RECT 69.500 46.195 69.760 46.620 ;
        RECT 70.000 45.180 70.230 46.415 ;
        RECT 70.790 45.180 71.020 46.415 ;
        RECT 71.380 45.180 71.610 46.415 ;
        RECT 61.980 43.810 62.240 44.600 ;
        RECT 58.840 43.580 60.080 43.810 ;
        RECT 61.000 43.580 62.240 43.810 ;
        RECT 64.175 43.810 64.435 44.690 ;
        RECT 64.675 43.970 64.905 44.860 ;
        RECT 65.465 43.970 65.695 44.860 ;
        RECT 66.055 43.970 66.285 44.860 ;
        RECT 66.845 43.970 67.075 44.935 ;
        RECT 69.985 44.860 70.245 45.180 ;
        RECT 70.775 44.860 71.035 45.180 ;
        RECT 71.365 44.860 71.625 45.180 ;
        RECT 72.170 45.105 72.400 46.415 ;
        RECT 72.590 45.545 72.850 46.620 ;
        RECT 73.010 45.105 73.180 47.045 ;
        RECT 72.170 44.935 73.180 45.105 ;
        RECT 73.325 44.935 73.680 47.045 ;
        RECT 74.060 47.320 74.415 49.515 ;
        RECT 75.335 49.450 75.565 50.415 ;
        RECT 76.125 49.540 76.355 50.415 ;
        RECT 76.715 49.540 76.945 50.415 ;
        RECT 77.505 49.540 77.735 50.415 ;
        RECT 77.975 49.785 78.235 50.575 ;
        RECT 80.160 50.575 81.400 50.805 ;
        RECT 82.320 50.575 83.560 50.805 ;
        RECT 80.160 49.880 80.420 50.575 ;
        RECT 74.555 49.280 75.565 49.450 ;
        RECT 74.555 47.320 74.725 49.280 ;
        RECT 74.885 47.765 75.145 48.900 ;
        RECT 75.335 47.970 75.565 49.280 ;
        RECT 76.110 49.220 76.370 49.540 ;
        RECT 76.700 49.220 76.960 49.540 ;
        RECT 77.490 49.220 77.750 49.540 ;
        RECT 76.125 47.970 76.355 49.220 ;
        RECT 76.715 47.970 76.945 49.220 ;
        RECT 77.505 47.970 77.735 49.220 ;
        RECT 77.975 47.765 78.235 48.270 ;
        RECT 74.885 47.535 76.075 47.765 ;
        RECT 76.995 47.535 78.235 47.765 ;
        RECT 78.660 47.320 79.015 49.510 ;
        RECT 74.060 47.045 74.725 47.320 ;
        RECT 78.345 47.045 79.015 47.320 ;
        RECT 74.060 44.940 74.415 47.045 ;
        RECT 74.835 46.620 76.075 46.850 ;
        RECT 76.995 46.620 78.185 46.850 ;
        RECT 74.835 46.195 75.095 46.620 ;
        RECT 75.335 45.180 75.565 46.415 ;
        RECT 76.125 45.180 76.355 46.415 ;
        RECT 76.715 45.180 76.945 46.415 ;
        RECT 67.315 43.810 67.575 44.600 ;
        RECT 64.175 43.580 65.415 43.810 ;
        RECT 66.335 43.580 67.575 43.810 ;
        RECT 69.500 43.810 69.760 44.690 ;
        RECT 70.000 43.970 70.230 44.860 ;
        RECT 70.790 43.970 71.020 44.860 ;
        RECT 71.380 43.970 71.610 44.860 ;
        RECT 72.170 43.970 72.400 44.935 ;
        RECT 75.320 44.860 75.580 45.180 ;
        RECT 76.110 44.860 76.370 45.180 ;
        RECT 76.700 44.860 76.960 45.180 ;
        RECT 77.505 45.105 77.735 46.415 ;
        RECT 77.925 45.545 78.185 46.620 ;
        RECT 78.345 45.105 78.515 47.045 ;
        RECT 77.505 44.935 78.515 45.105 ;
        RECT 78.660 44.935 79.015 47.045 ;
        RECT 79.385 47.320 79.740 49.515 ;
        RECT 80.660 49.450 80.890 50.415 ;
        RECT 81.450 49.540 81.680 50.415 ;
        RECT 82.040 49.540 82.270 50.415 ;
        RECT 82.830 49.540 83.060 50.415 ;
        RECT 83.300 49.785 83.560 50.575 ;
        RECT 85.495 50.575 86.735 50.805 ;
        RECT 87.655 50.575 88.895 50.805 ;
        RECT 85.495 49.880 85.755 50.575 ;
        RECT 79.880 49.280 80.890 49.450 ;
        RECT 79.880 47.320 80.050 49.280 ;
        RECT 80.210 47.765 80.470 48.900 ;
        RECT 80.660 47.970 80.890 49.280 ;
        RECT 81.435 49.220 81.695 49.540 ;
        RECT 82.025 49.220 82.285 49.540 ;
        RECT 82.815 49.220 83.075 49.540 ;
        RECT 81.450 47.970 81.680 49.220 ;
        RECT 82.040 47.970 82.270 49.220 ;
        RECT 82.830 47.970 83.060 49.220 ;
        RECT 83.300 47.765 83.560 48.270 ;
        RECT 80.210 47.535 81.400 47.765 ;
        RECT 82.320 47.535 83.560 47.765 ;
        RECT 83.985 47.320 84.340 49.510 ;
        RECT 79.385 47.045 80.050 47.320 ;
        RECT 83.670 47.045 84.340 47.320 ;
        RECT 79.385 44.940 79.740 47.045 ;
        RECT 80.160 46.620 81.400 46.850 ;
        RECT 82.320 46.620 83.510 46.850 ;
        RECT 80.160 46.195 80.420 46.620 ;
        RECT 80.660 45.180 80.890 46.415 ;
        RECT 81.450 45.180 81.680 46.415 ;
        RECT 82.040 45.180 82.270 46.415 ;
        RECT 72.640 43.810 72.900 44.600 ;
        RECT 69.500 43.580 70.740 43.810 ;
        RECT 71.660 43.580 72.900 43.810 ;
        RECT 74.835 43.810 75.095 44.690 ;
        RECT 75.335 43.970 75.565 44.860 ;
        RECT 76.125 43.970 76.355 44.860 ;
        RECT 76.715 43.970 76.945 44.860 ;
        RECT 77.505 43.970 77.735 44.935 ;
        RECT 80.645 44.860 80.905 45.180 ;
        RECT 81.435 44.860 81.695 45.180 ;
        RECT 82.025 44.860 82.285 45.180 ;
        RECT 82.830 45.105 83.060 46.415 ;
        RECT 83.250 45.545 83.510 46.620 ;
        RECT 83.670 45.105 83.840 47.045 ;
        RECT 82.830 44.935 83.840 45.105 ;
        RECT 83.985 44.935 84.340 47.045 ;
        RECT 84.720 47.320 85.075 49.515 ;
        RECT 85.995 49.450 86.225 50.415 ;
        RECT 86.785 49.540 87.015 50.415 ;
        RECT 87.375 49.540 87.605 50.415 ;
        RECT 88.165 49.540 88.395 50.415 ;
        RECT 88.635 49.785 88.895 50.575 ;
        RECT 90.820 50.575 92.060 50.805 ;
        RECT 92.980 50.575 94.220 50.805 ;
        RECT 90.820 49.880 91.080 50.575 ;
        RECT 85.215 49.280 86.225 49.450 ;
        RECT 85.215 47.320 85.385 49.280 ;
        RECT 85.545 47.765 85.805 48.900 ;
        RECT 85.995 47.970 86.225 49.280 ;
        RECT 86.770 49.220 87.030 49.540 ;
        RECT 87.360 49.220 87.620 49.540 ;
        RECT 88.150 49.220 88.410 49.540 ;
        RECT 86.785 47.970 87.015 49.220 ;
        RECT 87.375 47.970 87.605 49.220 ;
        RECT 88.165 47.970 88.395 49.220 ;
        RECT 88.635 47.765 88.895 48.270 ;
        RECT 85.545 47.535 86.735 47.765 ;
        RECT 87.655 47.535 88.895 47.765 ;
        RECT 89.320 47.320 89.675 49.510 ;
        RECT 84.720 47.045 85.385 47.320 ;
        RECT 89.005 47.045 89.675 47.320 ;
        RECT 84.720 44.940 85.075 47.045 ;
        RECT 85.495 46.620 86.735 46.850 ;
        RECT 87.655 46.620 88.845 46.850 ;
        RECT 85.495 46.195 85.755 46.620 ;
        RECT 85.995 45.180 86.225 46.415 ;
        RECT 86.785 45.180 87.015 46.415 ;
        RECT 87.375 45.180 87.605 46.415 ;
        RECT 77.975 43.810 78.235 44.600 ;
        RECT 74.835 43.580 76.075 43.810 ;
        RECT 76.995 43.580 78.235 43.810 ;
        RECT 80.160 43.810 80.420 44.690 ;
        RECT 80.660 43.970 80.890 44.860 ;
        RECT 81.450 43.970 81.680 44.860 ;
        RECT 82.040 43.970 82.270 44.860 ;
        RECT 82.830 43.970 83.060 44.935 ;
        RECT 85.980 44.860 86.240 45.180 ;
        RECT 86.770 44.860 87.030 45.180 ;
        RECT 87.360 44.860 87.620 45.180 ;
        RECT 88.165 45.105 88.395 46.415 ;
        RECT 88.585 45.545 88.845 46.620 ;
        RECT 89.005 45.105 89.175 47.045 ;
        RECT 88.165 44.935 89.175 45.105 ;
        RECT 89.320 44.935 89.675 47.045 ;
        RECT 90.045 47.320 90.400 49.515 ;
        RECT 91.320 49.450 91.550 50.415 ;
        RECT 92.110 49.540 92.340 50.415 ;
        RECT 92.700 49.540 92.930 50.415 ;
        RECT 93.490 49.540 93.720 50.415 ;
        RECT 93.960 49.785 94.220 50.575 ;
        RECT 96.155 50.575 97.395 50.805 ;
        RECT 98.315 50.575 99.555 50.805 ;
        RECT 96.155 49.880 96.415 50.575 ;
        RECT 90.540 49.280 91.550 49.450 ;
        RECT 90.540 47.320 90.710 49.280 ;
        RECT 90.870 47.765 91.130 48.900 ;
        RECT 91.320 47.970 91.550 49.280 ;
        RECT 92.095 49.220 92.355 49.540 ;
        RECT 92.685 49.220 92.945 49.540 ;
        RECT 93.475 49.220 93.735 49.540 ;
        RECT 92.110 47.970 92.340 49.220 ;
        RECT 92.700 47.970 92.930 49.220 ;
        RECT 93.490 47.970 93.720 49.220 ;
        RECT 93.960 47.765 94.220 48.270 ;
        RECT 90.870 47.535 92.060 47.765 ;
        RECT 92.980 47.535 94.220 47.765 ;
        RECT 94.645 47.320 95.000 49.510 ;
        RECT 90.045 47.045 90.710 47.320 ;
        RECT 94.330 47.045 95.000 47.320 ;
        RECT 90.045 44.940 90.400 47.045 ;
        RECT 90.820 46.620 92.060 46.850 ;
        RECT 92.980 46.620 94.170 46.850 ;
        RECT 90.820 46.195 91.080 46.620 ;
        RECT 91.320 45.180 91.550 46.415 ;
        RECT 92.110 45.180 92.340 46.415 ;
        RECT 92.700 45.180 92.930 46.415 ;
        RECT 83.300 43.810 83.560 44.600 ;
        RECT 80.160 43.580 81.400 43.810 ;
        RECT 82.320 43.580 83.560 43.810 ;
        RECT 85.495 43.810 85.755 44.690 ;
        RECT 85.995 43.970 86.225 44.860 ;
        RECT 86.785 43.970 87.015 44.860 ;
        RECT 87.375 43.970 87.605 44.860 ;
        RECT 88.165 43.970 88.395 44.935 ;
        RECT 91.305 44.860 91.565 45.180 ;
        RECT 92.095 44.860 92.355 45.180 ;
        RECT 92.685 44.860 92.945 45.180 ;
        RECT 93.490 45.105 93.720 46.415 ;
        RECT 93.910 45.545 94.170 46.620 ;
        RECT 94.330 45.105 94.500 47.045 ;
        RECT 93.490 44.935 94.500 45.105 ;
        RECT 94.645 44.935 95.000 47.045 ;
        RECT 95.380 47.320 95.735 49.515 ;
        RECT 96.655 49.450 96.885 50.415 ;
        RECT 97.445 49.540 97.675 50.415 ;
        RECT 98.035 49.540 98.265 50.415 ;
        RECT 98.825 49.540 99.055 50.415 ;
        RECT 99.295 49.785 99.555 50.575 ;
        RECT 101.480 50.575 102.720 50.805 ;
        RECT 103.640 50.575 104.880 50.805 ;
        RECT 101.480 49.880 101.740 50.575 ;
        RECT 95.875 49.280 96.885 49.450 ;
        RECT 95.875 47.320 96.045 49.280 ;
        RECT 96.205 47.765 96.465 48.900 ;
        RECT 96.655 47.970 96.885 49.280 ;
        RECT 97.430 49.220 97.690 49.540 ;
        RECT 98.020 49.220 98.280 49.540 ;
        RECT 98.810 49.220 99.070 49.540 ;
        RECT 97.445 47.970 97.675 49.220 ;
        RECT 98.035 47.970 98.265 49.220 ;
        RECT 98.825 47.970 99.055 49.220 ;
        RECT 99.295 47.765 99.555 48.270 ;
        RECT 96.205 47.535 97.395 47.765 ;
        RECT 98.315 47.535 99.555 47.765 ;
        RECT 99.980 47.320 100.335 49.510 ;
        RECT 95.380 47.045 96.045 47.320 ;
        RECT 99.665 47.045 100.335 47.320 ;
        RECT 95.380 44.940 95.735 47.045 ;
        RECT 96.155 46.620 97.395 46.850 ;
        RECT 98.315 46.620 99.505 46.850 ;
        RECT 96.155 46.195 96.415 46.620 ;
        RECT 96.655 45.180 96.885 46.415 ;
        RECT 97.445 45.180 97.675 46.415 ;
        RECT 98.035 45.180 98.265 46.415 ;
        RECT 88.635 43.810 88.895 44.600 ;
        RECT 85.495 43.580 86.735 43.810 ;
        RECT 87.655 43.580 88.895 43.810 ;
        RECT 90.820 43.810 91.080 44.690 ;
        RECT 91.320 43.970 91.550 44.860 ;
        RECT 92.110 43.970 92.340 44.860 ;
        RECT 92.700 43.970 92.930 44.860 ;
        RECT 93.490 43.970 93.720 44.935 ;
        RECT 96.640 44.860 96.900 45.180 ;
        RECT 97.430 44.860 97.690 45.180 ;
        RECT 98.020 44.860 98.280 45.180 ;
        RECT 98.825 45.105 99.055 46.415 ;
        RECT 99.245 45.545 99.505 46.620 ;
        RECT 99.665 45.105 99.835 47.045 ;
        RECT 98.825 44.935 99.835 45.105 ;
        RECT 99.980 44.935 100.335 47.045 ;
        RECT 100.705 47.320 101.060 49.515 ;
        RECT 101.980 49.450 102.210 50.415 ;
        RECT 102.770 49.540 103.000 50.415 ;
        RECT 103.360 49.540 103.590 50.415 ;
        RECT 104.150 49.540 104.380 50.415 ;
        RECT 104.620 49.785 104.880 50.575 ;
        RECT 106.815 50.575 108.055 50.805 ;
        RECT 108.975 50.575 110.215 50.805 ;
        RECT 106.815 49.880 107.075 50.575 ;
        RECT 101.200 49.280 102.210 49.450 ;
        RECT 101.200 47.320 101.370 49.280 ;
        RECT 101.530 47.765 101.790 48.900 ;
        RECT 101.980 47.970 102.210 49.280 ;
        RECT 102.755 49.220 103.015 49.540 ;
        RECT 103.345 49.220 103.605 49.540 ;
        RECT 104.135 49.220 104.395 49.540 ;
        RECT 102.770 47.970 103.000 49.220 ;
        RECT 103.360 47.970 103.590 49.220 ;
        RECT 104.150 47.970 104.380 49.220 ;
        RECT 104.620 47.765 104.880 48.270 ;
        RECT 101.530 47.535 102.720 47.765 ;
        RECT 103.640 47.535 104.880 47.765 ;
        RECT 105.305 47.320 105.660 49.510 ;
        RECT 100.705 47.045 101.370 47.320 ;
        RECT 104.990 47.045 105.660 47.320 ;
        RECT 100.705 44.940 101.060 47.045 ;
        RECT 101.480 46.620 102.720 46.850 ;
        RECT 103.640 46.620 104.830 46.850 ;
        RECT 101.480 46.195 101.740 46.620 ;
        RECT 101.980 45.180 102.210 46.415 ;
        RECT 102.770 45.180 103.000 46.415 ;
        RECT 103.360 45.180 103.590 46.415 ;
        RECT 93.960 43.810 94.220 44.600 ;
        RECT 90.820 43.580 92.060 43.810 ;
        RECT 92.980 43.580 94.220 43.810 ;
        RECT 96.155 43.810 96.415 44.690 ;
        RECT 96.655 43.970 96.885 44.860 ;
        RECT 97.445 43.970 97.675 44.860 ;
        RECT 98.035 43.970 98.265 44.860 ;
        RECT 98.825 43.970 99.055 44.935 ;
        RECT 101.965 44.860 102.225 45.180 ;
        RECT 102.755 44.860 103.015 45.180 ;
        RECT 103.345 44.860 103.605 45.180 ;
        RECT 104.150 45.105 104.380 46.415 ;
        RECT 104.570 45.545 104.830 46.620 ;
        RECT 104.990 45.105 105.160 47.045 ;
        RECT 104.150 44.935 105.160 45.105 ;
        RECT 105.305 44.935 105.660 47.045 ;
        RECT 106.040 47.320 106.395 49.515 ;
        RECT 107.315 49.450 107.545 50.415 ;
        RECT 108.105 49.540 108.335 50.415 ;
        RECT 108.695 49.540 108.925 50.415 ;
        RECT 109.485 49.540 109.715 50.415 ;
        RECT 109.955 49.785 110.215 50.575 ;
        RECT 112.140 50.575 113.380 50.805 ;
        RECT 114.300 50.575 115.540 50.805 ;
        RECT 112.140 49.880 112.400 50.575 ;
        RECT 106.535 49.280 107.545 49.450 ;
        RECT 106.535 47.320 106.705 49.280 ;
        RECT 106.865 47.765 107.125 48.900 ;
        RECT 107.315 47.970 107.545 49.280 ;
        RECT 108.090 49.220 108.350 49.540 ;
        RECT 108.680 49.220 108.940 49.540 ;
        RECT 109.470 49.220 109.730 49.540 ;
        RECT 108.105 47.970 108.335 49.220 ;
        RECT 108.695 47.970 108.925 49.220 ;
        RECT 109.485 47.970 109.715 49.220 ;
        RECT 109.955 47.765 110.215 48.270 ;
        RECT 106.865 47.535 108.055 47.765 ;
        RECT 108.975 47.535 110.215 47.765 ;
        RECT 110.640 47.320 110.995 49.510 ;
        RECT 106.040 47.045 106.705 47.320 ;
        RECT 110.325 47.045 110.995 47.320 ;
        RECT 106.040 44.940 106.395 47.045 ;
        RECT 106.815 46.620 108.055 46.850 ;
        RECT 108.975 46.620 110.165 46.850 ;
        RECT 106.815 46.195 107.075 46.620 ;
        RECT 107.315 45.180 107.545 46.415 ;
        RECT 108.105 45.180 108.335 46.415 ;
        RECT 108.695 45.180 108.925 46.415 ;
        RECT 99.295 43.810 99.555 44.600 ;
        RECT 96.155 43.580 97.395 43.810 ;
        RECT 98.315 43.580 99.555 43.810 ;
        RECT 101.480 43.810 101.740 44.690 ;
        RECT 101.980 43.970 102.210 44.860 ;
        RECT 102.770 43.970 103.000 44.860 ;
        RECT 103.360 43.970 103.590 44.860 ;
        RECT 104.150 43.970 104.380 44.935 ;
        RECT 107.300 44.860 107.560 45.180 ;
        RECT 108.090 44.860 108.350 45.180 ;
        RECT 108.680 44.860 108.940 45.180 ;
        RECT 109.485 45.105 109.715 46.415 ;
        RECT 109.905 45.545 110.165 46.620 ;
        RECT 110.325 45.105 110.495 47.045 ;
        RECT 109.485 44.935 110.495 45.105 ;
        RECT 110.640 44.935 110.995 47.045 ;
        RECT 111.365 47.320 111.720 49.515 ;
        RECT 112.640 49.450 112.870 50.415 ;
        RECT 113.430 49.540 113.660 50.415 ;
        RECT 114.020 49.540 114.250 50.415 ;
        RECT 114.810 49.540 115.040 50.415 ;
        RECT 115.280 49.785 115.540 50.575 ;
        RECT 117.475 50.575 118.715 50.805 ;
        RECT 119.635 50.575 120.875 50.805 ;
        RECT 117.475 49.880 117.735 50.575 ;
        RECT 111.860 49.280 112.870 49.450 ;
        RECT 111.860 47.320 112.030 49.280 ;
        RECT 112.190 47.765 112.450 48.900 ;
        RECT 112.640 47.970 112.870 49.280 ;
        RECT 113.415 49.220 113.675 49.540 ;
        RECT 114.005 49.220 114.265 49.540 ;
        RECT 114.795 49.220 115.055 49.540 ;
        RECT 113.430 47.970 113.660 49.220 ;
        RECT 114.020 47.970 114.250 49.220 ;
        RECT 114.810 47.970 115.040 49.220 ;
        RECT 115.280 47.765 115.540 48.270 ;
        RECT 112.190 47.535 113.380 47.765 ;
        RECT 114.300 47.535 115.540 47.765 ;
        RECT 115.965 47.320 116.320 49.510 ;
        RECT 111.365 47.045 112.030 47.320 ;
        RECT 115.650 47.045 116.320 47.320 ;
        RECT 111.365 44.940 111.720 47.045 ;
        RECT 112.140 46.620 113.380 46.850 ;
        RECT 114.300 46.620 115.490 46.850 ;
        RECT 112.140 46.195 112.400 46.620 ;
        RECT 112.640 45.180 112.870 46.415 ;
        RECT 113.430 45.180 113.660 46.415 ;
        RECT 114.020 45.180 114.250 46.415 ;
        RECT 104.620 43.810 104.880 44.600 ;
        RECT 101.480 43.580 102.720 43.810 ;
        RECT 103.640 43.580 104.880 43.810 ;
        RECT 106.815 43.810 107.075 44.690 ;
        RECT 107.315 43.970 107.545 44.860 ;
        RECT 108.105 43.970 108.335 44.860 ;
        RECT 108.695 43.970 108.925 44.860 ;
        RECT 109.485 43.970 109.715 44.935 ;
        RECT 112.625 44.860 112.885 45.180 ;
        RECT 113.415 44.860 113.675 45.180 ;
        RECT 114.005 44.860 114.265 45.180 ;
        RECT 114.810 45.105 115.040 46.415 ;
        RECT 115.230 45.545 115.490 46.620 ;
        RECT 115.650 45.105 115.820 47.045 ;
        RECT 114.810 44.935 115.820 45.105 ;
        RECT 115.965 44.935 116.320 47.045 ;
        RECT 116.700 47.320 117.055 49.515 ;
        RECT 117.975 49.450 118.205 50.415 ;
        RECT 118.765 49.540 118.995 50.415 ;
        RECT 119.355 49.540 119.585 50.415 ;
        RECT 120.145 49.540 120.375 50.415 ;
        RECT 120.615 49.785 120.875 50.575 ;
        RECT 117.195 49.280 118.205 49.450 ;
        RECT 117.195 47.320 117.365 49.280 ;
        RECT 117.525 47.765 117.785 48.900 ;
        RECT 117.975 47.970 118.205 49.280 ;
        RECT 118.750 49.220 119.010 49.540 ;
        RECT 119.340 49.220 119.600 49.540 ;
        RECT 120.130 49.220 120.390 49.540 ;
        RECT 118.765 47.970 118.995 49.220 ;
        RECT 119.355 47.970 119.585 49.220 ;
        RECT 120.145 47.970 120.375 49.220 ;
        RECT 120.615 47.765 120.875 48.270 ;
        RECT 117.525 47.535 118.715 47.765 ;
        RECT 119.635 47.535 120.875 47.765 ;
        RECT 121.300 47.320 121.655 49.510 ;
        RECT 116.700 47.045 117.365 47.320 ;
        RECT 120.985 47.045 121.655 47.320 ;
        RECT 116.700 44.940 117.055 47.045 ;
        RECT 117.475 46.620 118.715 46.850 ;
        RECT 119.635 46.620 120.825 46.850 ;
        RECT 117.475 46.195 117.735 46.620 ;
        RECT 117.975 45.180 118.205 46.415 ;
        RECT 118.765 45.180 118.995 46.415 ;
        RECT 119.355 45.180 119.585 46.415 ;
        RECT 109.955 43.810 110.215 44.600 ;
        RECT 106.815 43.580 108.055 43.810 ;
        RECT 108.975 43.580 110.215 43.810 ;
        RECT 112.140 43.810 112.400 44.690 ;
        RECT 112.640 43.970 112.870 44.860 ;
        RECT 113.430 43.970 113.660 44.860 ;
        RECT 114.020 43.970 114.250 44.860 ;
        RECT 114.810 43.970 115.040 44.935 ;
        RECT 117.960 44.860 118.220 45.180 ;
        RECT 118.750 44.860 119.010 45.180 ;
        RECT 119.340 44.860 119.600 45.180 ;
        RECT 120.145 45.105 120.375 46.415 ;
        RECT 120.565 45.545 120.825 46.620 ;
        RECT 120.985 45.105 121.155 47.045 ;
        RECT 120.145 44.935 121.155 45.105 ;
        RECT 121.300 44.935 121.655 47.045 ;
        RECT 122.025 47.320 122.380 49.530 ;
        RECT 123.300 49.450 123.530 50.415 ;
        RECT 124.090 49.540 124.320 50.415 ;
        RECT 124.680 49.540 124.910 50.415 ;
        RECT 125.470 49.540 125.700 50.415 ;
        RECT 122.520 49.280 123.530 49.450 ;
        RECT 122.520 47.320 122.690 49.280 ;
        RECT 123.300 47.970 123.530 49.280 ;
        RECT 124.075 49.220 124.335 49.540 ;
        RECT 124.665 49.220 124.925 49.540 ;
        RECT 125.455 49.220 125.715 49.540 ;
        RECT 124.090 47.970 124.320 49.220 ;
        RECT 124.680 47.970 124.910 49.220 ;
        RECT 125.470 47.970 125.700 49.220 ;
        RECT 126.625 47.320 126.980 49.530 ;
        RECT 122.025 47.045 122.690 47.320 ;
        RECT 126.310 47.045 126.980 47.320 ;
        RECT 122.025 44.955 122.380 47.045 ;
        RECT 123.300 45.180 123.530 46.415 ;
        RECT 124.090 45.180 124.320 46.415 ;
        RECT 124.680 45.180 124.910 46.415 ;
        RECT 115.280 43.810 115.540 44.600 ;
        RECT 112.140 43.580 113.380 43.810 ;
        RECT 114.300 43.580 115.540 43.810 ;
        RECT 117.475 43.810 117.735 44.690 ;
        RECT 117.975 43.970 118.205 44.860 ;
        RECT 118.765 43.970 118.995 44.860 ;
        RECT 119.355 43.970 119.585 44.860 ;
        RECT 120.145 43.970 120.375 44.935 ;
        RECT 123.285 44.860 123.545 45.180 ;
        RECT 124.075 44.860 124.335 45.180 ;
        RECT 124.665 44.860 124.925 45.180 ;
        RECT 125.470 45.105 125.700 46.415 ;
        RECT 126.310 45.105 126.480 47.045 ;
        RECT 125.470 44.935 126.480 45.105 ;
        RECT 126.625 44.955 126.980 47.045 ;
        RECT 120.615 43.810 120.875 44.600 ;
        RECT 123.300 43.970 123.530 44.860 ;
        RECT 124.090 43.970 124.320 44.860 ;
        RECT 124.680 43.970 124.910 44.860 ;
        RECT 125.470 43.970 125.700 44.935 ;
        RECT 117.475 43.580 118.715 43.810 ;
        RECT 119.635 43.580 120.875 43.810 ;
        RECT 12.425 43.240 12.715 43.255 ;
        RECT 37.520 43.040 38.760 43.270 ;
        RECT 39.680 43.040 40.920 43.270 ;
        RECT 10.510 39.735 10.810 41.185 ;
        RECT 15.985 41.020 25.285 41.255 ;
        RECT 11.745 40.635 13.345 40.925 ;
        RECT 14.165 40.635 20.945 40.870 ;
        RECT 16.040 40.450 17.645 40.480 ;
        RECT 21.425 40.450 25.285 41.020 ;
        RECT 15.985 40.255 25.285 40.450 ;
        RECT 15.985 40.215 25.710 40.255 ;
        RECT 16.040 40.190 17.645 40.215 ;
        RECT 23.850 39.215 25.710 40.215 ;
        RECT 31.420 39.785 31.775 41.995 ;
        RECT 32.695 41.915 32.925 42.880 ;
        RECT 33.485 42.005 33.715 42.880 ;
        RECT 34.075 42.005 34.305 42.880 ;
        RECT 34.865 42.005 35.095 42.880 ;
        RECT 37.520 42.345 37.780 43.040 ;
        RECT 31.915 41.745 32.925 41.915 ;
        RECT 31.915 39.785 32.085 41.745 ;
        RECT 32.695 40.435 32.925 41.745 ;
        RECT 33.470 41.685 33.730 42.005 ;
        RECT 34.060 41.685 34.320 42.005 ;
        RECT 34.850 41.685 35.110 42.005 ;
        RECT 33.485 40.435 33.715 41.685 ;
        RECT 34.075 40.435 34.305 41.685 ;
        RECT 34.865 40.435 35.095 41.685 ;
        RECT 36.020 39.785 36.375 41.995 ;
        RECT 31.420 39.510 32.085 39.785 ;
        RECT 35.705 39.510 36.375 39.785 ;
        RECT 31.420 37.420 31.775 39.510 ;
        RECT 32.695 37.645 32.925 38.880 ;
        RECT 33.485 37.645 33.715 38.880 ;
        RECT 34.075 37.645 34.305 38.880 ;
        RECT 32.680 37.325 32.940 37.645 ;
        RECT 33.470 37.325 33.730 37.645 ;
        RECT 34.060 37.325 34.320 37.645 ;
        RECT 34.865 37.570 35.095 38.880 ;
        RECT 35.705 37.570 35.875 39.510 ;
        RECT 34.865 37.400 35.875 37.570 ;
        RECT 36.020 37.420 36.375 39.510 ;
        RECT 36.745 39.785 37.100 41.980 ;
        RECT 38.020 41.915 38.250 42.880 ;
        RECT 38.810 42.005 39.040 42.880 ;
        RECT 39.400 42.005 39.630 42.880 ;
        RECT 40.190 42.005 40.420 42.880 ;
        RECT 40.660 42.250 40.920 43.040 ;
        RECT 42.855 43.040 44.095 43.270 ;
        RECT 45.015 43.040 46.255 43.270 ;
        RECT 42.855 42.345 43.115 43.040 ;
        RECT 37.240 41.745 38.250 41.915 ;
        RECT 37.240 39.785 37.410 41.745 ;
        RECT 37.570 40.230 37.830 41.365 ;
        RECT 38.020 40.435 38.250 41.745 ;
        RECT 38.795 41.685 39.055 42.005 ;
        RECT 39.385 41.685 39.645 42.005 ;
        RECT 40.175 41.685 40.435 42.005 ;
        RECT 38.810 40.435 39.040 41.685 ;
        RECT 39.400 40.435 39.630 41.685 ;
        RECT 40.190 40.435 40.420 41.685 ;
        RECT 40.660 40.230 40.920 40.735 ;
        RECT 37.570 40.000 38.760 40.230 ;
        RECT 39.680 40.000 40.920 40.230 ;
        RECT 41.345 39.785 41.700 41.975 ;
        RECT 36.745 39.510 37.410 39.785 ;
        RECT 41.030 39.510 41.700 39.785 ;
        RECT 36.745 37.405 37.100 39.510 ;
        RECT 37.520 39.085 38.760 39.315 ;
        RECT 39.680 39.085 40.870 39.315 ;
        RECT 37.520 38.660 37.780 39.085 ;
        RECT 38.020 37.645 38.250 38.880 ;
        RECT 38.810 37.645 39.040 38.880 ;
        RECT 39.400 37.645 39.630 38.880 ;
        RECT 10.500 36.190 10.820 36.675 ;
        RECT 16.115 36.300 25.305 36.535 ;
        RECT 32.695 36.435 32.925 37.325 ;
        RECT 33.485 36.435 33.715 37.325 ;
        RECT 34.075 36.435 34.305 37.325 ;
        RECT 34.865 36.435 35.095 37.400 ;
        RECT 38.005 37.325 38.265 37.645 ;
        RECT 38.795 37.325 39.055 37.645 ;
        RECT 39.385 37.325 39.645 37.645 ;
        RECT 40.190 37.570 40.420 38.880 ;
        RECT 40.610 38.010 40.870 39.085 ;
        RECT 41.030 37.570 41.200 39.510 ;
        RECT 40.190 37.400 41.200 37.570 ;
        RECT 41.345 37.400 41.700 39.510 ;
        RECT 42.080 39.785 42.435 41.980 ;
        RECT 43.355 41.915 43.585 42.880 ;
        RECT 44.145 42.005 44.375 42.880 ;
        RECT 44.735 42.005 44.965 42.880 ;
        RECT 45.525 42.005 45.755 42.880 ;
        RECT 45.995 42.250 46.255 43.040 ;
        RECT 48.180 43.040 49.420 43.270 ;
        RECT 50.340 43.040 51.580 43.270 ;
        RECT 48.180 42.345 48.440 43.040 ;
        RECT 42.575 41.745 43.585 41.915 ;
        RECT 42.575 39.785 42.745 41.745 ;
        RECT 42.905 40.230 43.165 41.365 ;
        RECT 43.355 40.435 43.585 41.745 ;
        RECT 44.130 41.685 44.390 42.005 ;
        RECT 44.720 41.685 44.980 42.005 ;
        RECT 45.510 41.685 45.770 42.005 ;
        RECT 44.145 40.435 44.375 41.685 ;
        RECT 44.735 40.435 44.965 41.685 ;
        RECT 45.525 40.435 45.755 41.685 ;
        RECT 45.995 40.230 46.255 40.735 ;
        RECT 42.905 40.000 44.095 40.230 ;
        RECT 45.015 40.000 46.255 40.230 ;
        RECT 46.680 39.785 47.035 41.975 ;
        RECT 42.080 39.510 42.745 39.785 ;
        RECT 46.365 39.510 47.035 39.785 ;
        RECT 42.080 37.405 42.435 39.510 ;
        RECT 42.855 39.085 44.095 39.315 ;
        RECT 45.015 39.085 46.205 39.315 ;
        RECT 42.855 38.660 43.115 39.085 ;
        RECT 43.355 37.645 43.585 38.880 ;
        RECT 44.145 37.645 44.375 38.880 ;
        RECT 44.735 37.645 44.965 38.880 ;
        RECT 10.500 35.860 11.960 36.190 ;
        RECT 10.500 35.640 10.820 35.860 ;
        RECT 12.400 35.115 12.720 36.105 ;
        RECT 14.585 35.860 16.005 36.185 ;
        RECT 19.990 35.730 25.305 36.300 ;
        RECT 37.520 36.275 37.780 37.155 ;
        RECT 38.020 36.435 38.250 37.325 ;
        RECT 38.810 36.435 39.040 37.325 ;
        RECT 39.400 36.435 39.630 37.325 ;
        RECT 40.190 36.435 40.420 37.400 ;
        RECT 43.340 37.325 43.600 37.645 ;
        RECT 44.130 37.325 44.390 37.645 ;
        RECT 44.720 37.325 44.980 37.645 ;
        RECT 45.525 37.570 45.755 38.880 ;
        RECT 45.945 38.010 46.205 39.085 ;
        RECT 46.365 37.570 46.535 39.510 ;
        RECT 45.525 37.400 46.535 37.570 ;
        RECT 46.680 37.400 47.035 39.510 ;
        RECT 47.405 39.785 47.760 41.980 ;
        RECT 48.680 41.915 48.910 42.880 ;
        RECT 49.470 42.005 49.700 42.880 ;
        RECT 50.060 42.005 50.290 42.880 ;
        RECT 50.850 42.005 51.080 42.880 ;
        RECT 51.320 42.250 51.580 43.040 ;
        RECT 53.515 43.040 54.755 43.270 ;
        RECT 55.675 43.040 56.915 43.270 ;
        RECT 53.515 42.345 53.775 43.040 ;
        RECT 47.900 41.745 48.910 41.915 ;
        RECT 47.900 39.785 48.070 41.745 ;
        RECT 48.230 40.230 48.490 41.365 ;
        RECT 48.680 40.435 48.910 41.745 ;
        RECT 49.455 41.685 49.715 42.005 ;
        RECT 50.045 41.685 50.305 42.005 ;
        RECT 50.835 41.685 51.095 42.005 ;
        RECT 49.470 40.435 49.700 41.685 ;
        RECT 50.060 40.435 50.290 41.685 ;
        RECT 50.850 40.435 51.080 41.685 ;
        RECT 51.320 40.230 51.580 40.735 ;
        RECT 48.230 40.000 49.420 40.230 ;
        RECT 50.340 40.000 51.580 40.230 ;
        RECT 52.005 39.785 52.360 41.975 ;
        RECT 47.405 39.510 48.070 39.785 ;
        RECT 51.690 39.510 52.360 39.785 ;
        RECT 47.405 37.405 47.760 39.510 ;
        RECT 48.180 39.085 49.420 39.315 ;
        RECT 50.340 39.085 51.530 39.315 ;
        RECT 48.180 38.660 48.440 39.085 ;
        RECT 48.680 37.645 48.910 38.880 ;
        RECT 49.470 37.645 49.700 38.880 ;
        RECT 50.060 37.645 50.290 38.880 ;
        RECT 40.660 36.275 40.920 37.065 ;
        RECT 37.520 36.045 38.760 36.275 ;
        RECT 39.680 36.045 40.920 36.275 ;
        RECT 42.855 36.275 43.115 37.155 ;
        RECT 43.355 36.435 43.585 37.325 ;
        RECT 44.145 36.435 44.375 37.325 ;
        RECT 44.735 36.435 44.965 37.325 ;
        RECT 45.525 36.435 45.755 37.400 ;
        RECT 48.665 37.325 48.925 37.645 ;
        RECT 49.455 37.325 49.715 37.645 ;
        RECT 50.045 37.325 50.305 37.645 ;
        RECT 50.850 37.570 51.080 38.880 ;
        RECT 51.270 38.010 51.530 39.085 ;
        RECT 51.690 37.570 51.860 39.510 ;
        RECT 50.850 37.400 51.860 37.570 ;
        RECT 52.005 37.400 52.360 39.510 ;
        RECT 52.740 39.785 53.095 41.980 ;
        RECT 54.015 41.915 54.245 42.880 ;
        RECT 54.805 42.005 55.035 42.880 ;
        RECT 55.395 42.005 55.625 42.880 ;
        RECT 56.185 42.005 56.415 42.880 ;
        RECT 56.655 42.250 56.915 43.040 ;
        RECT 58.840 43.040 60.080 43.270 ;
        RECT 61.000 43.040 62.240 43.270 ;
        RECT 58.840 42.345 59.100 43.040 ;
        RECT 53.235 41.745 54.245 41.915 ;
        RECT 53.235 39.785 53.405 41.745 ;
        RECT 53.565 40.230 53.825 41.365 ;
        RECT 54.015 40.435 54.245 41.745 ;
        RECT 54.790 41.685 55.050 42.005 ;
        RECT 55.380 41.685 55.640 42.005 ;
        RECT 56.170 41.685 56.430 42.005 ;
        RECT 54.805 40.435 55.035 41.685 ;
        RECT 55.395 40.435 55.625 41.685 ;
        RECT 56.185 40.435 56.415 41.685 ;
        RECT 56.655 40.230 56.915 40.735 ;
        RECT 53.565 40.000 54.755 40.230 ;
        RECT 55.675 40.000 56.915 40.230 ;
        RECT 57.340 39.785 57.695 41.975 ;
        RECT 52.740 39.510 53.405 39.785 ;
        RECT 57.025 39.510 57.695 39.785 ;
        RECT 52.740 37.405 53.095 39.510 ;
        RECT 53.515 39.085 54.755 39.315 ;
        RECT 55.675 39.085 56.865 39.315 ;
        RECT 53.515 38.660 53.775 39.085 ;
        RECT 54.015 37.645 54.245 38.880 ;
        RECT 54.805 37.645 55.035 38.880 ;
        RECT 55.395 37.645 55.625 38.880 ;
        RECT 45.995 36.275 46.255 37.065 ;
        RECT 42.855 36.045 44.095 36.275 ;
        RECT 45.015 36.045 46.255 36.275 ;
        RECT 48.180 36.275 48.440 37.155 ;
        RECT 48.680 36.435 48.910 37.325 ;
        RECT 49.470 36.435 49.700 37.325 ;
        RECT 50.060 36.435 50.290 37.325 ;
        RECT 50.850 36.435 51.080 37.400 ;
        RECT 54.000 37.325 54.260 37.645 ;
        RECT 54.790 37.325 55.050 37.645 ;
        RECT 55.380 37.325 55.640 37.645 ;
        RECT 56.185 37.570 56.415 38.880 ;
        RECT 56.605 38.010 56.865 39.085 ;
        RECT 57.025 37.570 57.195 39.510 ;
        RECT 56.185 37.400 57.195 37.570 ;
        RECT 57.340 37.400 57.695 39.510 ;
        RECT 58.065 39.785 58.420 41.980 ;
        RECT 59.340 41.915 59.570 42.880 ;
        RECT 60.130 42.005 60.360 42.880 ;
        RECT 60.720 42.005 60.950 42.880 ;
        RECT 61.510 42.005 61.740 42.880 ;
        RECT 61.980 42.250 62.240 43.040 ;
        RECT 64.175 43.040 65.415 43.270 ;
        RECT 66.335 43.040 67.575 43.270 ;
        RECT 64.175 42.345 64.435 43.040 ;
        RECT 58.560 41.745 59.570 41.915 ;
        RECT 58.560 39.785 58.730 41.745 ;
        RECT 58.890 40.230 59.150 41.365 ;
        RECT 59.340 40.435 59.570 41.745 ;
        RECT 60.115 41.685 60.375 42.005 ;
        RECT 60.705 41.685 60.965 42.005 ;
        RECT 61.495 41.685 61.755 42.005 ;
        RECT 60.130 40.435 60.360 41.685 ;
        RECT 60.720 40.435 60.950 41.685 ;
        RECT 61.510 40.435 61.740 41.685 ;
        RECT 61.980 40.230 62.240 40.735 ;
        RECT 58.890 40.000 60.080 40.230 ;
        RECT 61.000 40.000 62.240 40.230 ;
        RECT 62.665 39.785 63.020 41.975 ;
        RECT 58.065 39.510 58.730 39.785 ;
        RECT 62.350 39.510 63.020 39.785 ;
        RECT 58.065 37.405 58.420 39.510 ;
        RECT 58.840 39.085 60.080 39.315 ;
        RECT 61.000 39.085 62.190 39.315 ;
        RECT 58.840 38.660 59.100 39.085 ;
        RECT 59.340 37.645 59.570 38.880 ;
        RECT 60.130 37.645 60.360 38.880 ;
        RECT 60.720 37.645 60.950 38.880 ;
        RECT 51.320 36.275 51.580 37.065 ;
        RECT 48.180 36.045 49.420 36.275 ;
        RECT 50.340 36.045 51.580 36.275 ;
        RECT 53.515 36.275 53.775 37.155 ;
        RECT 54.015 36.435 54.245 37.325 ;
        RECT 54.805 36.435 55.035 37.325 ;
        RECT 55.395 36.435 55.625 37.325 ;
        RECT 56.185 36.435 56.415 37.400 ;
        RECT 59.325 37.325 59.585 37.645 ;
        RECT 60.115 37.325 60.375 37.645 ;
        RECT 60.705 37.325 60.965 37.645 ;
        RECT 61.510 37.570 61.740 38.880 ;
        RECT 61.930 38.010 62.190 39.085 ;
        RECT 62.350 37.570 62.520 39.510 ;
        RECT 61.510 37.400 62.520 37.570 ;
        RECT 62.665 37.400 63.020 39.510 ;
        RECT 63.400 39.785 63.755 41.980 ;
        RECT 64.675 41.915 64.905 42.880 ;
        RECT 65.465 42.005 65.695 42.880 ;
        RECT 66.055 42.005 66.285 42.880 ;
        RECT 66.845 42.005 67.075 42.880 ;
        RECT 67.315 42.250 67.575 43.040 ;
        RECT 69.500 43.040 70.740 43.270 ;
        RECT 71.660 43.040 72.900 43.270 ;
        RECT 69.500 42.345 69.760 43.040 ;
        RECT 63.895 41.745 64.905 41.915 ;
        RECT 63.895 39.785 64.065 41.745 ;
        RECT 64.225 40.230 64.485 41.365 ;
        RECT 64.675 40.435 64.905 41.745 ;
        RECT 65.450 41.685 65.710 42.005 ;
        RECT 66.040 41.685 66.300 42.005 ;
        RECT 66.830 41.685 67.090 42.005 ;
        RECT 65.465 40.435 65.695 41.685 ;
        RECT 66.055 40.435 66.285 41.685 ;
        RECT 66.845 40.435 67.075 41.685 ;
        RECT 67.315 40.230 67.575 40.735 ;
        RECT 64.225 40.000 65.415 40.230 ;
        RECT 66.335 40.000 67.575 40.230 ;
        RECT 68.000 39.785 68.355 41.975 ;
        RECT 63.400 39.510 64.065 39.785 ;
        RECT 67.685 39.510 68.355 39.785 ;
        RECT 63.400 37.405 63.755 39.510 ;
        RECT 64.175 39.085 65.415 39.315 ;
        RECT 66.335 39.085 67.525 39.315 ;
        RECT 64.175 38.660 64.435 39.085 ;
        RECT 64.675 37.645 64.905 38.880 ;
        RECT 65.465 37.645 65.695 38.880 ;
        RECT 66.055 37.645 66.285 38.880 ;
        RECT 56.655 36.275 56.915 37.065 ;
        RECT 53.515 36.045 54.755 36.275 ;
        RECT 55.675 36.045 56.915 36.275 ;
        RECT 58.840 36.275 59.100 37.155 ;
        RECT 59.340 36.435 59.570 37.325 ;
        RECT 60.130 36.435 60.360 37.325 ;
        RECT 60.720 36.435 60.950 37.325 ;
        RECT 61.510 36.435 61.740 37.400 ;
        RECT 64.660 37.325 64.920 37.645 ;
        RECT 65.450 37.325 65.710 37.645 ;
        RECT 66.040 37.325 66.300 37.645 ;
        RECT 66.845 37.570 67.075 38.880 ;
        RECT 67.265 38.010 67.525 39.085 ;
        RECT 67.685 37.570 67.855 39.510 ;
        RECT 66.845 37.400 67.855 37.570 ;
        RECT 68.000 37.400 68.355 39.510 ;
        RECT 68.725 39.785 69.080 41.980 ;
        RECT 70.000 41.915 70.230 42.880 ;
        RECT 70.790 42.005 71.020 42.880 ;
        RECT 71.380 42.005 71.610 42.880 ;
        RECT 72.170 42.005 72.400 42.880 ;
        RECT 72.640 42.250 72.900 43.040 ;
        RECT 74.835 43.040 76.075 43.270 ;
        RECT 76.995 43.040 78.235 43.270 ;
        RECT 74.835 42.345 75.095 43.040 ;
        RECT 69.220 41.745 70.230 41.915 ;
        RECT 69.220 39.785 69.390 41.745 ;
        RECT 69.550 40.230 69.810 41.365 ;
        RECT 70.000 40.435 70.230 41.745 ;
        RECT 70.775 41.685 71.035 42.005 ;
        RECT 71.365 41.685 71.625 42.005 ;
        RECT 72.155 41.685 72.415 42.005 ;
        RECT 70.790 40.435 71.020 41.685 ;
        RECT 71.380 40.435 71.610 41.685 ;
        RECT 72.170 40.435 72.400 41.685 ;
        RECT 72.640 40.230 72.900 40.735 ;
        RECT 69.550 40.000 70.740 40.230 ;
        RECT 71.660 40.000 72.900 40.230 ;
        RECT 73.325 39.785 73.680 41.975 ;
        RECT 68.725 39.510 69.390 39.785 ;
        RECT 73.010 39.510 73.680 39.785 ;
        RECT 68.725 37.405 69.080 39.510 ;
        RECT 69.500 39.085 70.740 39.315 ;
        RECT 71.660 39.085 72.850 39.315 ;
        RECT 69.500 38.660 69.760 39.085 ;
        RECT 70.000 37.645 70.230 38.880 ;
        RECT 70.790 37.645 71.020 38.880 ;
        RECT 71.380 37.645 71.610 38.880 ;
        RECT 61.980 36.275 62.240 37.065 ;
        RECT 58.840 36.045 60.080 36.275 ;
        RECT 61.000 36.045 62.240 36.275 ;
        RECT 64.175 36.275 64.435 37.155 ;
        RECT 64.675 36.435 64.905 37.325 ;
        RECT 65.465 36.435 65.695 37.325 ;
        RECT 66.055 36.435 66.285 37.325 ;
        RECT 66.845 36.435 67.075 37.400 ;
        RECT 69.985 37.325 70.245 37.645 ;
        RECT 70.775 37.325 71.035 37.645 ;
        RECT 71.365 37.325 71.625 37.645 ;
        RECT 72.170 37.570 72.400 38.880 ;
        RECT 72.590 38.010 72.850 39.085 ;
        RECT 73.010 37.570 73.180 39.510 ;
        RECT 72.170 37.400 73.180 37.570 ;
        RECT 73.325 37.400 73.680 39.510 ;
        RECT 74.060 39.785 74.415 41.980 ;
        RECT 75.335 41.915 75.565 42.880 ;
        RECT 76.125 42.005 76.355 42.880 ;
        RECT 76.715 42.005 76.945 42.880 ;
        RECT 77.505 42.005 77.735 42.880 ;
        RECT 77.975 42.250 78.235 43.040 ;
        RECT 80.160 43.040 81.400 43.270 ;
        RECT 82.320 43.040 83.560 43.270 ;
        RECT 80.160 42.345 80.420 43.040 ;
        RECT 74.555 41.745 75.565 41.915 ;
        RECT 74.555 39.785 74.725 41.745 ;
        RECT 74.885 40.230 75.145 41.365 ;
        RECT 75.335 40.435 75.565 41.745 ;
        RECT 76.110 41.685 76.370 42.005 ;
        RECT 76.700 41.685 76.960 42.005 ;
        RECT 77.490 41.685 77.750 42.005 ;
        RECT 76.125 40.435 76.355 41.685 ;
        RECT 76.715 40.435 76.945 41.685 ;
        RECT 77.505 40.435 77.735 41.685 ;
        RECT 77.975 40.230 78.235 40.735 ;
        RECT 74.885 40.000 76.075 40.230 ;
        RECT 76.995 40.000 78.235 40.230 ;
        RECT 78.660 39.785 79.015 41.975 ;
        RECT 74.060 39.510 74.725 39.785 ;
        RECT 78.345 39.510 79.015 39.785 ;
        RECT 74.060 37.405 74.415 39.510 ;
        RECT 74.835 39.085 76.075 39.315 ;
        RECT 76.995 39.085 78.185 39.315 ;
        RECT 74.835 38.660 75.095 39.085 ;
        RECT 75.335 37.645 75.565 38.880 ;
        RECT 76.125 37.645 76.355 38.880 ;
        RECT 76.715 37.645 76.945 38.880 ;
        RECT 67.315 36.275 67.575 37.065 ;
        RECT 64.175 36.045 65.415 36.275 ;
        RECT 66.335 36.045 67.575 36.275 ;
        RECT 69.500 36.275 69.760 37.155 ;
        RECT 70.000 36.435 70.230 37.325 ;
        RECT 70.790 36.435 71.020 37.325 ;
        RECT 71.380 36.435 71.610 37.325 ;
        RECT 72.170 36.435 72.400 37.400 ;
        RECT 75.320 37.325 75.580 37.645 ;
        RECT 76.110 37.325 76.370 37.645 ;
        RECT 76.700 37.325 76.960 37.645 ;
        RECT 77.505 37.570 77.735 38.880 ;
        RECT 77.925 38.010 78.185 39.085 ;
        RECT 78.345 37.570 78.515 39.510 ;
        RECT 77.505 37.400 78.515 37.570 ;
        RECT 78.660 37.400 79.015 39.510 ;
        RECT 79.385 39.785 79.740 41.980 ;
        RECT 80.660 41.915 80.890 42.880 ;
        RECT 81.450 42.005 81.680 42.880 ;
        RECT 82.040 42.005 82.270 42.880 ;
        RECT 82.830 42.005 83.060 42.880 ;
        RECT 83.300 42.250 83.560 43.040 ;
        RECT 85.495 43.040 86.735 43.270 ;
        RECT 87.655 43.040 88.895 43.270 ;
        RECT 85.495 42.345 85.755 43.040 ;
        RECT 79.880 41.745 80.890 41.915 ;
        RECT 79.880 39.785 80.050 41.745 ;
        RECT 80.210 40.230 80.470 41.365 ;
        RECT 80.660 40.435 80.890 41.745 ;
        RECT 81.435 41.685 81.695 42.005 ;
        RECT 82.025 41.685 82.285 42.005 ;
        RECT 82.815 41.685 83.075 42.005 ;
        RECT 81.450 40.435 81.680 41.685 ;
        RECT 82.040 40.435 82.270 41.685 ;
        RECT 82.830 40.435 83.060 41.685 ;
        RECT 83.300 40.230 83.560 40.735 ;
        RECT 80.210 40.000 81.400 40.230 ;
        RECT 82.320 40.000 83.560 40.230 ;
        RECT 83.985 39.785 84.340 41.975 ;
        RECT 79.385 39.510 80.050 39.785 ;
        RECT 83.670 39.510 84.340 39.785 ;
        RECT 79.385 37.405 79.740 39.510 ;
        RECT 80.160 39.085 81.400 39.315 ;
        RECT 82.320 39.085 83.510 39.315 ;
        RECT 80.160 38.660 80.420 39.085 ;
        RECT 80.660 37.645 80.890 38.880 ;
        RECT 81.450 37.645 81.680 38.880 ;
        RECT 82.040 37.645 82.270 38.880 ;
        RECT 72.640 36.275 72.900 37.065 ;
        RECT 69.500 36.045 70.740 36.275 ;
        RECT 71.660 36.045 72.900 36.275 ;
        RECT 74.835 36.275 75.095 37.155 ;
        RECT 75.335 36.435 75.565 37.325 ;
        RECT 76.125 36.435 76.355 37.325 ;
        RECT 76.715 36.435 76.945 37.325 ;
        RECT 77.505 36.435 77.735 37.400 ;
        RECT 80.645 37.325 80.905 37.645 ;
        RECT 81.435 37.325 81.695 37.645 ;
        RECT 82.025 37.325 82.285 37.645 ;
        RECT 82.830 37.570 83.060 38.880 ;
        RECT 83.250 38.010 83.510 39.085 ;
        RECT 83.670 37.570 83.840 39.510 ;
        RECT 82.830 37.400 83.840 37.570 ;
        RECT 83.985 37.400 84.340 39.510 ;
        RECT 84.720 39.785 85.075 41.980 ;
        RECT 85.995 41.915 86.225 42.880 ;
        RECT 86.785 42.005 87.015 42.880 ;
        RECT 87.375 42.005 87.605 42.880 ;
        RECT 88.165 42.005 88.395 42.880 ;
        RECT 88.635 42.250 88.895 43.040 ;
        RECT 90.820 43.040 92.060 43.270 ;
        RECT 92.980 43.040 94.220 43.270 ;
        RECT 90.820 42.345 91.080 43.040 ;
        RECT 85.215 41.745 86.225 41.915 ;
        RECT 85.215 39.785 85.385 41.745 ;
        RECT 85.545 40.230 85.805 41.365 ;
        RECT 85.995 40.435 86.225 41.745 ;
        RECT 86.770 41.685 87.030 42.005 ;
        RECT 87.360 41.685 87.620 42.005 ;
        RECT 88.150 41.685 88.410 42.005 ;
        RECT 86.785 40.435 87.015 41.685 ;
        RECT 87.375 40.435 87.605 41.685 ;
        RECT 88.165 40.435 88.395 41.685 ;
        RECT 88.635 40.230 88.895 40.735 ;
        RECT 85.545 40.000 86.735 40.230 ;
        RECT 87.655 40.000 88.895 40.230 ;
        RECT 89.320 39.785 89.675 41.975 ;
        RECT 84.720 39.510 85.385 39.785 ;
        RECT 89.005 39.510 89.675 39.785 ;
        RECT 84.720 37.405 85.075 39.510 ;
        RECT 85.495 39.085 86.735 39.315 ;
        RECT 87.655 39.085 88.845 39.315 ;
        RECT 85.495 38.660 85.755 39.085 ;
        RECT 85.995 37.645 86.225 38.880 ;
        RECT 86.785 37.645 87.015 38.880 ;
        RECT 87.375 37.645 87.605 38.880 ;
        RECT 77.975 36.275 78.235 37.065 ;
        RECT 74.835 36.045 76.075 36.275 ;
        RECT 76.995 36.045 78.235 36.275 ;
        RECT 80.160 36.275 80.420 37.155 ;
        RECT 80.660 36.435 80.890 37.325 ;
        RECT 81.450 36.435 81.680 37.325 ;
        RECT 82.040 36.435 82.270 37.325 ;
        RECT 82.830 36.435 83.060 37.400 ;
        RECT 85.980 37.325 86.240 37.645 ;
        RECT 86.770 37.325 87.030 37.645 ;
        RECT 87.360 37.325 87.620 37.645 ;
        RECT 88.165 37.570 88.395 38.880 ;
        RECT 88.585 38.010 88.845 39.085 ;
        RECT 89.005 37.570 89.175 39.510 ;
        RECT 88.165 37.400 89.175 37.570 ;
        RECT 89.320 37.400 89.675 39.510 ;
        RECT 90.045 39.785 90.400 41.980 ;
        RECT 91.320 41.915 91.550 42.880 ;
        RECT 92.110 42.005 92.340 42.880 ;
        RECT 92.700 42.005 92.930 42.880 ;
        RECT 93.490 42.005 93.720 42.880 ;
        RECT 93.960 42.250 94.220 43.040 ;
        RECT 96.155 43.040 97.395 43.270 ;
        RECT 98.315 43.040 99.555 43.270 ;
        RECT 96.155 42.345 96.415 43.040 ;
        RECT 90.540 41.745 91.550 41.915 ;
        RECT 90.540 39.785 90.710 41.745 ;
        RECT 90.870 40.230 91.130 41.365 ;
        RECT 91.320 40.435 91.550 41.745 ;
        RECT 92.095 41.685 92.355 42.005 ;
        RECT 92.685 41.685 92.945 42.005 ;
        RECT 93.475 41.685 93.735 42.005 ;
        RECT 92.110 40.435 92.340 41.685 ;
        RECT 92.700 40.435 92.930 41.685 ;
        RECT 93.490 40.435 93.720 41.685 ;
        RECT 93.960 40.230 94.220 40.735 ;
        RECT 90.870 40.000 92.060 40.230 ;
        RECT 92.980 40.000 94.220 40.230 ;
        RECT 94.645 39.785 95.000 41.975 ;
        RECT 90.045 39.510 90.710 39.785 ;
        RECT 94.330 39.510 95.000 39.785 ;
        RECT 90.045 37.405 90.400 39.510 ;
        RECT 90.820 39.085 92.060 39.315 ;
        RECT 92.980 39.085 94.170 39.315 ;
        RECT 90.820 38.660 91.080 39.085 ;
        RECT 91.320 37.645 91.550 38.880 ;
        RECT 92.110 37.645 92.340 38.880 ;
        RECT 92.700 37.645 92.930 38.880 ;
        RECT 83.300 36.275 83.560 37.065 ;
        RECT 80.160 36.045 81.400 36.275 ;
        RECT 82.320 36.045 83.560 36.275 ;
        RECT 85.495 36.275 85.755 37.155 ;
        RECT 85.995 36.435 86.225 37.325 ;
        RECT 86.785 36.435 87.015 37.325 ;
        RECT 87.375 36.435 87.605 37.325 ;
        RECT 88.165 36.435 88.395 37.400 ;
        RECT 91.305 37.325 91.565 37.645 ;
        RECT 92.095 37.325 92.355 37.645 ;
        RECT 92.685 37.325 92.945 37.645 ;
        RECT 93.490 37.570 93.720 38.880 ;
        RECT 93.910 38.010 94.170 39.085 ;
        RECT 94.330 37.570 94.500 39.510 ;
        RECT 93.490 37.400 94.500 37.570 ;
        RECT 94.645 37.400 95.000 39.510 ;
        RECT 95.380 39.785 95.735 41.980 ;
        RECT 96.655 41.915 96.885 42.880 ;
        RECT 97.445 42.005 97.675 42.880 ;
        RECT 98.035 42.005 98.265 42.880 ;
        RECT 98.825 42.005 99.055 42.880 ;
        RECT 99.295 42.250 99.555 43.040 ;
        RECT 101.480 43.040 102.720 43.270 ;
        RECT 103.640 43.040 104.880 43.270 ;
        RECT 101.480 42.345 101.740 43.040 ;
        RECT 95.875 41.745 96.885 41.915 ;
        RECT 95.875 39.785 96.045 41.745 ;
        RECT 96.205 40.230 96.465 41.365 ;
        RECT 96.655 40.435 96.885 41.745 ;
        RECT 97.430 41.685 97.690 42.005 ;
        RECT 98.020 41.685 98.280 42.005 ;
        RECT 98.810 41.685 99.070 42.005 ;
        RECT 97.445 40.435 97.675 41.685 ;
        RECT 98.035 40.435 98.265 41.685 ;
        RECT 98.825 40.435 99.055 41.685 ;
        RECT 99.295 40.230 99.555 40.735 ;
        RECT 96.205 40.000 97.395 40.230 ;
        RECT 98.315 40.000 99.555 40.230 ;
        RECT 99.980 39.785 100.335 41.975 ;
        RECT 95.380 39.510 96.045 39.785 ;
        RECT 99.665 39.510 100.335 39.785 ;
        RECT 95.380 37.405 95.735 39.510 ;
        RECT 96.155 39.085 97.395 39.315 ;
        RECT 98.315 39.085 99.505 39.315 ;
        RECT 96.155 38.660 96.415 39.085 ;
        RECT 96.655 37.645 96.885 38.880 ;
        RECT 97.445 37.645 97.675 38.880 ;
        RECT 98.035 37.645 98.265 38.880 ;
        RECT 88.635 36.275 88.895 37.065 ;
        RECT 85.495 36.045 86.735 36.275 ;
        RECT 87.655 36.045 88.895 36.275 ;
        RECT 90.820 36.275 91.080 37.155 ;
        RECT 91.320 36.435 91.550 37.325 ;
        RECT 92.110 36.435 92.340 37.325 ;
        RECT 92.700 36.435 92.930 37.325 ;
        RECT 93.490 36.435 93.720 37.400 ;
        RECT 96.640 37.325 96.900 37.645 ;
        RECT 97.430 37.325 97.690 37.645 ;
        RECT 98.020 37.325 98.280 37.645 ;
        RECT 98.825 37.570 99.055 38.880 ;
        RECT 99.245 38.010 99.505 39.085 ;
        RECT 99.665 37.570 99.835 39.510 ;
        RECT 98.825 37.400 99.835 37.570 ;
        RECT 99.980 37.400 100.335 39.510 ;
        RECT 100.705 39.785 101.060 41.980 ;
        RECT 101.980 41.915 102.210 42.880 ;
        RECT 102.770 42.005 103.000 42.880 ;
        RECT 103.360 42.005 103.590 42.880 ;
        RECT 104.150 42.005 104.380 42.880 ;
        RECT 104.620 42.250 104.880 43.040 ;
        RECT 106.815 43.040 108.055 43.270 ;
        RECT 108.975 43.040 110.215 43.270 ;
        RECT 106.815 42.345 107.075 43.040 ;
        RECT 101.200 41.745 102.210 41.915 ;
        RECT 101.200 39.785 101.370 41.745 ;
        RECT 101.530 40.230 101.790 41.365 ;
        RECT 101.980 40.435 102.210 41.745 ;
        RECT 102.755 41.685 103.015 42.005 ;
        RECT 103.345 41.685 103.605 42.005 ;
        RECT 104.135 41.685 104.395 42.005 ;
        RECT 102.770 40.435 103.000 41.685 ;
        RECT 103.360 40.435 103.590 41.685 ;
        RECT 104.150 40.435 104.380 41.685 ;
        RECT 104.620 40.230 104.880 40.735 ;
        RECT 101.530 40.000 102.720 40.230 ;
        RECT 103.640 40.000 104.880 40.230 ;
        RECT 105.305 39.785 105.660 41.975 ;
        RECT 100.705 39.510 101.370 39.785 ;
        RECT 104.990 39.510 105.660 39.785 ;
        RECT 100.705 37.405 101.060 39.510 ;
        RECT 101.480 39.085 102.720 39.315 ;
        RECT 103.640 39.085 104.830 39.315 ;
        RECT 101.480 38.660 101.740 39.085 ;
        RECT 101.980 37.645 102.210 38.880 ;
        RECT 102.770 37.645 103.000 38.880 ;
        RECT 103.360 37.645 103.590 38.880 ;
        RECT 93.960 36.275 94.220 37.065 ;
        RECT 90.820 36.045 92.060 36.275 ;
        RECT 92.980 36.045 94.220 36.275 ;
        RECT 96.155 36.275 96.415 37.155 ;
        RECT 96.655 36.435 96.885 37.325 ;
        RECT 97.445 36.435 97.675 37.325 ;
        RECT 98.035 36.435 98.265 37.325 ;
        RECT 98.825 36.435 99.055 37.400 ;
        RECT 101.965 37.325 102.225 37.645 ;
        RECT 102.755 37.325 103.015 37.645 ;
        RECT 103.345 37.325 103.605 37.645 ;
        RECT 104.150 37.570 104.380 38.880 ;
        RECT 104.570 38.010 104.830 39.085 ;
        RECT 104.990 37.570 105.160 39.510 ;
        RECT 104.150 37.400 105.160 37.570 ;
        RECT 105.305 37.400 105.660 39.510 ;
        RECT 106.040 39.785 106.395 41.980 ;
        RECT 107.315 41.915 107.545 42.880 ;
        RECT 108.105 42.005 108.335 42.880 ;
        RECT 108.695 42.005 108.925 42.880 ;
        RECT 109.485 42.005 109.715 42.880 ;
        RECT 109.955 42.250 110.215 43.040 ;
        RECT 112.140 43.040 113.380 43.270 ;
        RECT 114.300 43.040 115.540 43.270 ;
        RECT 112.140 42.345 112.400 43.040 ;
        RECT 106.535 41.745 107.545 41.915 ;
        RECT 106.535 39.785 106.705 41.745 ;
        RECT 106.865 40.230 107.125 41.365 ;
        RECT 107.315 40.435 107.545 41.745 ;
        RECT 108.090 41.685 108.350 42.005 ;
        RECT 108.680 41.685 108.940 42.005 ;
        RECT 109.470 41.685 109.730 42.005 ;
        RECT 108.105 40.435 108.335 41.685 ;
        RECT 108.695 40.435 108.925 41.685 ;
        RECT 109.485 40.435 109.715 41.685 ;
        RECT 109.955 40.230 110.215 40.735 ;
        RECT 106.865 40.000 108.055 40.230 ;
        RECT 108.975 40.000 110.215 40.230 ;
        RECT 110.640 39.785 110.995 41.975 ;
        RECT 106.040 39.510 106.705 39.785 ;
        RECT 110.325 39.510 110.995 39.785 ;
        RECT 106.040 37.405 106.395 39.510 ;
        RECT 106.815 39.085 108.055 39.315 ;
        RECT 108.975 39.085 110.165 39.315 ;
        RECT 106.815 38.660 107.075 39.085 ;
        RECT 107.315 37.645 107.545 38.880 ;
        RECT 108.105 37.645 108.335 38.880 ;
        RECT 108.695 37.645 108.925 38.880 ;
        RECT 99.295 36.275 99.555 37.065 ;
        RECT 96.155 36.045 97.395 36.275 ;
        RECT 98.315 36.045 99.555 36.275 ;
        RECT 101.480 36.275 101.740 37.155 ;
        RECT 101.980 36.435 102.210 37.325 ;
        RECT 102.770 36.435 103.000 37.325 ;
        RECT 103.360 36.435 103.590 37.325 ;
        RECT 104.150 36.435 104.380 37.400 ;
        RECT 107.300 37.325 107.560 37.645 ;
        RECT 108.090 37.325 108.350 37.645 ;
        RECT 108.680 37.325 108.940 37.645 ;
        RECT 109.485 37.570 109.715 38.880 ;
        RECT 109.905 38.010 110.165 39.085 ;
        RECT 110.325 37.570 110.495 39.510 ;
        RECT 109.485 37.400 110.495 37.570 ;
        RECT 110.640 37.400 110.995 39.510 ;
        RECT 111.365 39.785 111.720 41.980 ;
        RECT 112.640 41.915 112.870 42.880 ;
        RECT 113.430 42.005 113.660 42.880 ;
        RECT 114.020 42.005 114.250 42.880 ;
        RECT 114.810 42.005 115.040 42.880 ;
        RECT 115.280 42.250 115.540 43.040 ;
        RECT 117.475 43.040 118.715 43.270 ;
        RECT 119.635 43.040 120.875 43.270 ;
        RECT 117.475 42.345 117.735 43.040 ;
        RECT 111.860 41.745 112.870 41.915 ;
        RECT 111.860 39.785 112.030 41.745 ;
        RECT 112.190 40.230 112.450 41.365 ;
        RECT 112.640 40.435 112.870 41.745 ;
        RECT 113.415 41.685 113.675 42.005 ;
        RECT 114.005 41.685 114.265 42.005 ;
        RECT 114.795 41.685 115.055 42.005 ;
        RECT 113.430 40.435 113.660 41.685 ;
        RECT 114.020 40.435 114.250 41.685 ;
        RECT 114.810 40.435 115.040 41.685 ;
        RECT 115.280 40.230 115.540 40.735 ;
        RECT 112.190 40.000 113.380 40.230 ;
        RECT 114.300 40.000 115.540 40.230 ;
        RECT 115.965 39.785 116.320 41.975 ;
        RECT 111.365 39.510 112.030 39.785 ;
        RECT 115.650 39.510 116.320 39.785 ;
        RECT 111.365 37.405 111.720 39.510 ;
        RECT 112.140 39.085 113.380 39.315 ;
        RECT 114.300 39.085 115.490 39.315 ;
        RECT 112.140 38.660 112.400 39.085 ;
        RECT 112.640 37.645 112.870 38.880 ;
        RECT 113.430 37.645 113.660 38.880 ;
        RECT 114.020 37.645 114.250 38.880 ;
        RECT 104.620 36.275 104.880 37.065 ;
        RECT 101.480 36.045 102.720 36.275 ;
        RECT 103.640 36.045 104.880 36.275 ;
        RECT 106.815 36.275 107.075 37.155 ;
        RECT 107.315 36.435 107.545 37.325 ;
        RECT 108.105 36.435 108.335 37.325 ;
        RECT 108.695 36.435 108.925 37.325 ;
        RECT 109.485 36.435 109.715 37.400 ;
        RECT 112.625 37.325 112.885 37.645 ;
        RECT 113.415 37.325 113.675 37.645 ;
        RECT 114.005 37.325 114.265 37.645 ;
        RECT 114.810 37.570 115.040 38.880 ;
        RECT 115.230 38.010 115.490 39.085 ;
        RECT 115.650 37.570 115.820 39.510 ;
        RECT 114.810 37.400 115.820 37.570 ;
        RECT 115.965 37.400 116.320 39.510 ;
        RECT 116.700 39.785 117.055 41.980 ;
        RECT 117.975 41.915 118.205 42.880 ;
        RECT 118.765 42.005 118.995 42.880 ;
        RECT 119.355 42.005 119.585 42.880 ;
        RECT 120.145 42.005 120.375 42.880 ;
        RECT 120.615 42.250 120.875 43.040 ;
        RECT 117.195 41.745 118.205 41.915 ;
        RECT 117.195 39.785 117.365 41.745 ;
        RECT 117.525 40.230 117.785 41.365 ;
        RECT 117.975 40.435 118.205 41.745 ;
        RECT 118.750 41.685 119.010 42.005 ;
        RECT 119.340 41.685 119.600 42.005 ;
        RECT 120.130 41.685 120.390 42.005 ;
        RECT 118.765 40.435 118.995 41.685 ;
        RECT 119.355 40.435 119.585 41.685 ;
        RECT 120.145 40.435 120.375 41.685 ;
        RECT 120.615 40.230 120.875 40.735 ;
        RECT 117.525 40.000 118.715 40.230 ;
        RECT 119.635 40.000 120.875 40.230 ;
        RECT 121.300 39.785 121.655 41.975 ;
        RECT 116.700 39.510 117.365 39.785 ;
        RECT 120.985 39.510 121.655 39.785 ;
        RECT 116.700 37.405 117.055 39.510 ;
        RECT 117.475 39.085 118.715 39.315 ;
        RECT 119.635 39.085 120.825 39.315 ;
        RECT 117.475 38.660 117.735 39.085 ;
        RECT 117.975 37.645 118.205 38.880 ;
        RECT 118.765 37.645 118.995 38.880 ;
        RECT 119.355 37.645 119.585 38.880 ;
        RECT 109.955 36.275 110.215 37.065 ;
        RECT 106.815 36.045 108.055 36.275 ;
        RECT 108.975 36.045 110.215 36.275 ;
        RECT 112.140 36.275 112.400 37.155 ;
        RECT 112.640 36.435 112.870 37.325 ;
        RECT 113.430 36.435 113.660 37.325 ;
        RECT 114.020 36.435 114.250 37.325 ;
        RECT 114.810 36.435 115.040 37.400 ;
        RECT 117.960 37.325 118.220 37.645 ;
        RECT 118.750 37.325 119.010 37.645 ;
        RECT 119.340 37.325 119.600 37.645 ;
        RECT 120.145 37.570 120.375 38.880 ;
        RECT 120.565 38.010 120.825 39.085 ;
        RECT 120.985 37.570 121.155 39.510 ;
        RECT 120.145 37.400 121.155 37.570 ;
        RECT 121.300 37.400 121.655 39.510 ;
        RECT 122.025 39.785 122.380 41.995 ;
        RECT 123.300 41.915 123.530 42.880 ;
        RECT 124.090 42.005 124.320 42.880 ;
        RECT 124.680 42.005 124.910 42.880 ;
        RECT 125.470 42.005 125.700 42.880 ;
        RECT 122.520 41.745 123.530 41.915 ;
        RECT 122.520 39.785 122.690 41.745 ;
        RECT 123.300 40.435 123.530 41.745 ;
        RECT 124.075 41.685 124.335 42.005 ;
        RECT 124.665 41.685 124.925 42.005 ;
        RECT 125.455 41.685 125.715 42.005 ;
        RECT 124.090 40.435 124.320 41.685 ;
        RECT 124.680 40.435 124.910 41.685 ;
        RECT 125.470 40.435 125.700 41.685 ;
        RECT 126.625 39.785 126.980 41.995 ;
        RECT 122.025 39.510 122.690 39.785 ;
        RECT 126.310 39.510 126.980 39.785 ;
        RECT 122.025 37.420 122.380 39.510 ;
        RECT 123.300 37.645 123.530 38.880 ;
        RECT 124.090 37.645 124.320 38.880 ;
        RECT 124.680 37.645 124.910 38.880 ;
        RECT 115.280 36.275 115.540 37.065 ;
        RECT 112.140 36.045 113.380 36.275 ;
        RECT 114.300 36.045 115.540 36.275 ;
        RECT 117.475 36.275 117.735 37.155 ;
        RECT 117.975 36.435 118.205 37.325 ;
        RECT 118.765 36.435 118.995 37.325 ;
        RECT 119.355 36.435 119.585 37.325 ;
        RECT 120.145 36.435 120.375 37.400 ;
        RECT 123.285 37.325 123.545 37.645 ;
        RECT 124.075 37.325 124.335 37.645 ;
        RECT 124.665 37.325 124.925 37.645 ;
        RECT 125.470 37.570 125.700 38.880 ;
        RECT 126.310 37.570 126.480 39.510 ;
        RECT 125.470 37.400 126.480 37.570 ;
        RECT 126.625 37.420 126.980 39.510 ;
        RECT 120.615 36.275 120.875 37.065 ;
        RECT 123.300 36.435 123.530 37.325 ;
        RECT 124.090 36.435 124.320 37.325 ;
        RECT 124.680 36.435 124.910 37.325 ;
        RECT 125.470 36.435 125.700 37.400 ;
        RECT 117.475 36.045 118.715 36.275 ;
        RECT 119.635 36.045 120.875 36.275 ;
        RECT 16.115 35.495 25.305 35.730 ;
        RECT 37.520 35.505 38.760 35.735 ;
        RECT 39.680 35.505 40.920 35.735 ;
        RECT 12.425 35.100 12.715 35.115 ;
        RECT 26.145 33.115 26.405 33.120 ;
        RECT 10.510 31.595 10.810 33.045 ;
        RECT 15.985 32.880 26.455 33.115 ;
        RECT 11.745 32.495 13.345 32.785 ;
        RECT 14.165 32.495 20.945 32.730 ;
        RECT 16.040 32.310 17.645 32.340 ;
        RECT 21.425 32.310 26.455 32.880 ;
        RECT 15.985 32.075 26.455 32.310 ;
        RECT 31.420 32.250 31.775 34.460 ;
        RECT 32.695 34.380 32.925 35.345 ;
        RECT 33.485 34.470 33.715 35.345 ;
        RECT 34.075 34.470 34.305 35.345 ;
        RECT 34.865 34.470 35.095 35.345 ;
        RECT 37.520 34.810 37.780 35.505 ;
        RECT 31.915 34.210 32.925 34.380 ;
        RECT 31.915 32.250 32.085 34.210 ;
        RECT 32.695 32.900 32.925 34.210 ;
        RECT 33.470 34.150 33.730 34.470 ;
        RECT 34.060 34.150 34.320 34.470 ;
        RECT 34.850 34.150 35.110 34.470 ;
        RECT 33.485 32.900 33.715 34.150 ;
        RECT 34.075 32.900 34.305 34.150 ;
        RECT 34.865 32.900 35.095 34.150 ;
        RECT 36.020 32.250 36.375 34.460 ;
        RECT 16.040 32.050 17.645 32.075 ;
        RECT 31.420 31.975 32.085 32.250 ;
        RECT 35.705 31.975 36.375 32.250 ;
        RECT 31.420 29.885 31.775 31.975 ;
        RECT 32.695 30.110 32.925 31.345 ;
        RECT 33.485 30.110 33.715 31.345 ;
        RECT 34.075 30.110 34.305 31.345 ;
        RECT 32.680 29.790 32.940 30.110 ;
        RECT 33.470 29.790 33.730 30.110 ;
        RECT 34.060 29.790 34.320 30.110 ;
        RECT 34.865 30.035 35.095 31.345 ;
        RECT 35.705 30.035 35.875 31.975 ;
        RECT 34.865 29.865 35.875 30.035 ;
        RECT 36.020 29.885 36.375 31.975 ;
        RECT 36.745 32.250 37.100 34.445 ;
        RECT 38.020 34.380 38.250 35.345 ;
        RECT 38.810 34.470 39.040 35.345 ;
        RECT 39.400 34.470 39.630 35.345 ;
        RECT 40.190 34.470 40.420 35.345 ;
        RECT 40.660 34.715 40.920 35.505 ;
        RECT 42.855 35.505 44.095 35.735 ;
        RECT 45.015 35.505 46.255 35.735 ;
        RECT 42.855 34.810 43.115 35.505 ;
        RECT 37.240 34.210 38.250 34.380 ;
        RECT 37.240 32.250 37.410 34.210 ;
        RECT 37.570 32.695 37.830 33.830 ;
        RECT 38.020 32.900 38.250 34.210 ;
        RECT 38.795 34.150 39.055 34.470 ;
        RECT 39.385 34.150 39.645 34.470 ;
        RECT 40.175 34.150 40.435 34.470 ;
        RECT 38.810 32.900 39.040 34.150 ;
        RECT 39.400 32.900 39.630 34.150 ;
        RECT 40.190 32.900 40.420 34.150 ;
        RECT 40.660 32.695 40.920 33.200 ;
        RECT 37.570 32.465 38.760 32.695 ;
        RECT 39.680 32.465 40.920 32.695 ;
        RECT 41.345 32.250 41.700 34.440 ;
        RECT 36.745 31.975 37.410 32.250 ;
        RECT 41.030 31.975 41.700 32.250 ;
        RECT 36.745 29.870 37.100 31.975 ;
        RECT 37.520 31.550 38.760 31.780 ;
        RECT 39.680 31.550 40.870 31.780 ;
        RECT 37.520 31.125 37.780 31.550 ;
        RECT 38.020 30.110 38.250 31.345 ;
        RECT 38.810 30.110 39.040 31.345 ;
        RECT 39.400 30.110 39.630 31.345 ;
        RECT 32.695 28.900 32.925 29.790 ;
        RECT 33.485 28.900 33.715 29.790 ;
        RECT 34.075 28.900 34.305 29.790 ;
        RECT 34.865 28.900 35.095 29.865 ;
        RECT 38.005 29.790 38.265 30.110 ;
        RECT 38.795 29.790 39.055 30.110 ;
        RECT 39.385 29.790 39.645 30.110 ;
        RECT 40.190 30.035 40.420 31.345 ;
        RECT 40.610 30.475 40.870 31.550 ;
        RECT 41.030 30.035 41.200 31.975 ;
        RECT 40.190 29.865 41.200 30.035 ;
        RECT 41.345 29.865 41.700 31.975 ;
        RECT 42.080 32.250 42.435 34.445 ;
        RECT 43.355 34.380 43.585 35.345 ;
        RECT 44.145 34.470 44.375 35.345 ;
        RECT 44.735 34.470 44.965 35.345 ;
        RECT 45.525 34.470 45.755 35.345 ;
        RECT 45.995 34.715 46.255 35.505 ;
        RECT 48.180 35.505 49.420 35.735 ;
        RECT 50.340 35.505 51.580 35.735 ;
        RECT 48.180 34.810 48.440 35.505 ;
        RECT 42.575 34.210 43.585 34.380 ;
        RECT 42.575 32.250 42.745 34.210 ;
        RECT 42.905 32.695 43.165 33.830 ;
        RECT 43.355 32.900 43.585 34.210 ;
        RECT 44.130 34.150 44.390 34.470 ;
        RECT 44.720 34.150 44.980 34.470 ;
        RECT 45.510 34.150 45.770 34.470 ;
        RECT 44.145 32.900 44.375 34.150 ;
        RECT 44.735 32.900 44.965 34.150 ;
        RECT 45.525 32.900 45.755 34.150 ;
        RECT 45.995 32.695 46.255 33.200 ;
        RECT 42.905 32.465 44.095 32.695 ;
        RECT 45.015 32.465 46.255 32.695 ;
        RECT 46.680 32.250 47.035 34.440 ;
        RECT 42.080 31.975 42.745 32.250 ;
        RECT 46.365 31.975 47.035 32.250 ;
        RECT 42.080 29.870 42.435 31.975 ;
        RECT 42.855 31.550 44.095 31.780 ;
        RECT 45.015 31.550 46.205 31.780 ;
        RECT 42.855 31.125 43.115 31.550 ;
        RECT 43.355 30.110 43.585 31.345 ;
        RECT 44.145 30.110 44.375 31.345 ;
        RECT 44.735 30.110 44.965 31.345 ;
        RECT 37.520 28.740 37.780 29.620 ;
        RECT 38.020 28.900 38.250 29.790 ;
        RECT 38.810 28.900 39.040 29.790 ;
        RECT 39.400 28.900 39.630 29.790 ;
        RECT 40.190 28.900 40.420 29.865 ;
        RECT 43.340 29.790 43.600 30.110 ;
        RECT 44.130 29.790 44.390 30.110 ;
        RECT 44.720 29.790 44.980 30.110 ;
        RECT 45.525 30.035 45.755 31.345 ;
        RECT 45.945 30.475 46.205 31.550 ;
        RECT 46.365 30.035 46.535 31.975 ;
        RECT 45.525 29.865 46.535 30.035 ;
        RECT 46.680 29.865 47.035 31.975 ;
        RECT 47.405 32.250 47.760 34.445 ;
        RECT 48.680 34.380 48.910 35.345 ;
        RECT 49.470 34.470 49.700 35.345 ;
        RECT 50.060 34.470 50.290 35.345 ;
        RECT 50.850 34.470 51.080 35.345 ;
        RECT 51.320 34.715 51.580 35.505 ;
        RECT 53.515 35.505 54.755 35.735 ;
        RECT 55.675 35.505 56.915 35.735 ;
        RECT 53.515 34.810 53.775 35.505 ;
        RECT 47.900 34.210 48.910 34.380 ;
        RECT 47.900 32.250 48.070 34.210 ;
        RECT 48.230 32.695 48.490 33.830 ;
        RECT 48.680 32.900 48.910 34.210 ;
        RECT 49.455 34.150 49.715 34.470 ;
        RECT 50.045 34.150 50.305 34.470 ;
        RECT 50.835 34.150 51.095 34.470 ;
        RECT 49.470 32.900 49.700 34.150 ;
        RECT 50.060 32.900 50.290 34.150 ;
        RECT 50.850 32.900 51.080 34.150 ;
        RECT 51.320 32.695 51.580 33.200 ;
        RECT 48.230 32.465 49.420 32.695 ;
        RECT 50.340 32.465 51.580 32.695 ;
        RECT 52.005 32.250 52.360 34.440 ;
        RECT 47.405 31.975 48.070 32.250 ;
        RECT 51.690 31.975 52.360 32.250 ;
        RECT 47.405 29.870 47.760 31.975 ;
        RECT 48.180 31.550 49.420 31.780 ;
        RECT 50.340 31.550 51.530 31.780 ;
        RECT 48.180 31.125 48.440 31.550 ;
        RECT 48.680 30.110 48.910 31.345 ;
        RECT 49.470 30.110 49.700 31.345 ;
        RECT 50.060 30.110 50.290 31.345 ;
        RECT 40.660 28.740 40.920 29.530 ;
        RECT 10.500 28.050 10.820 28.535 ;
        RECT 37.520 28.510 38.760 28.740 ;
        RECT 39.680 28.510 40.920 28.740 ;
        RECT 42.855 28.740 43.115 29.620 ;
        RECT 43.355 28.900 43.585 29.790 ;
        RECT 44.145 28.900 44.375 29.790 ;
        RECT 44.735 28.900 44.965 29.790 ;
        RECT 45.525 28.900 45.755 29.865 ;
        RECT 48.665 29.790 48.925 30.110 ;
        RECT 49.455 29.790 49.715 30.110 ;
        RECT 50.045 29.790 50.305 30.110 ;
        RECT 50.850 30.035 51.080 31.345 ;
        RECT 51.270 30.475 51.530 31.550 ;
        RECT 51.690 30.035 51.860 31.975 ;
        RECT 50.850 29.865 51.860 30.035 ;
        RECT 52.005 29.865 52.360 31.975 ;
        RECT 52.740 32.250 53.095 34.445 ;
        RECT 54.015 34.380 54.245 35.345 ;
        RECT 54.805 34.470 55.035 35.345 ;
        RECT 55.395 34.470 55.625 35.345 ;
        RECT 56.185 34.470 56.415 35.345 ;
        RECT 56.655 34.715 56.915 35.505 ;
        RECT 58.840 35.505 60.080 35.735 ;
        RECT 61.000 35.505 62.240 35.735 ;
        RECT 58.840 34.810 59.100 35.505 ;
        RECT 53.235 34.210 54.245 34.380 ;
        RECT 53.235 32.250 53.405 34.210 ;
        RECT 53.565 32.695 53.825 33.830 ;
        RECT 54.015 32.900 54.245 34.210 ;
        RECT 54.790 34.150 55.050 34.470 ;
        RECT 55.380 34.150 55.640 34.470 ;
        RECT 56.170 34.150 56.430 34.470 ;
        RECT 54.805 32.900 55.035 34.150 ;
        RECT 55.395 32.900 55.625 34.150 ;
        RECT 56.185 32.900 56.415 34.150 ;
        RECT 56.655 32.695 56.915 33.200 ;
        RECT 53.565 32.465 54.755 32.695 ;
        RECT 55.675 32.465 56.915 32.695 ;
        RECT 57.340 32.250 57.695 34.440 ;
        RECT 52.740 31.975 53.405 32.250 ;
        RECT 57.025 31.975 57.695 32.250 ;
        RECT 52.740 29.870 53.095 31.975 ;
        RECT 53.515 31.550 54.755 31.780 ;
        RECT 55.675 31.550 56.865 31.780 ;
        RECT 53.515 31.125 53.775 31.550 ;
        RECT 54.015 30.110 54.245 31.345 ;
        RECT 54.805 30.110 55.035 31.345 ;
        RECT 55.395 30.110 55.625 31.345 ;
        RECT 45.995 28.740 46.255 29.530 ;
        RECT 42.855 28.510 44.095 28.740 ;
        RECT 45.015 28.510 46.255 28.740 ;
        RECT 48.180 28.740 48.440 29.620 ;
        RECT 48.680 28.900 48.910 29.790 ;
        RECT 49.470 28.900 49.700 29.790 ;
        RECT 50.060 28.900 50.290 29.790 ;
        RECT 50.850 28.900 51.080 29.865 ;
        RECT 54.000 29.790 54.260 30.110 ;
        RECT 54.790 29.790 55.050 30.110 ;
        RECT 55.380 29.790 55.640 30.110 ;
        RECT 56.185 30.035 56.415 31.345 ;
        RECT 56.605 30.475 56.865 31.550 ;
        RECT 57.025 30.035 57.195 31.975 ;
        RECT 56.185 29.865 57.195 30.035 ;
        RECT 57.340 29.865 57.695 31.975 ;
        RECT 58.065 32.250 58.420 34.445 ;
        RECT 59.340 34.380 59.570 35.345 ;
        RECT 60.130 34.470 60.360 35.345 ;
        RECT 60.720 34.470 60.950 35.345 ;
        RECT 61.510 34.470 61.740 35.345 ;
        RECT 61.980 34.715 62.240 35.505 ;
        RECT 64.175 35.505 65.415 35.735 ;
        RECT 66.335 35.505 67.575 35.735 ;
        RECT 64.175 34.810 64.435 35.505 ;
        RECT 58.560 34.210 59.570 34.380 ;
        RECT 58.560 32.250 58.730 34.210 ;
        RECT 58.890 32.695 59.150 33.830 ;
        RECT 59.340 32.900 59.570 34.210 ;
        RECT 60.115 34.150 60.375 34.470 ;
        RECT 60.705 34.150 60.965 34.470 ;
        RECT 61.495 34.150 61.755 34.470 ;
        RECT 60.130 32.900 60.360 34.150 ;
        RECT 60.720 32.900 60.950 34.150 ;
        RECT 61.510 32.900 61.740 34.150 ;
        RECT 61.980 32.695 62.240 33.200 ;
        RECT 58.890 32.465 60.080 32.695 ;
        RECT 61.000 32.465 62.240 32.695 ;
        RECT 62.665 32.250 63.020 34.440 ;
        RECT 58.065 31.975 58.730 32.250 ;
        RECT 62.350 31.975 63.020 32.250 ;
        RECT 58.065 29.870 58.420 31.975 ;
        RECT 58.840 31.550 60.080 31.780 ;
        RECT 61.000 31.550 62.190 31.780 ;
        RECT 58.840 31.125 59.100 31.550 ;
        RECT 59.340 30.110 59.570 31.345 ;
        RECT 60.130 30.110 60.360 31.345 ;
        RECT 60.720 30.110 60.950 31.345 ;
        RECT 51.320 28.740 51.580 29.530 ;
        RECT 48.180 28.510 49.420 28.740 ;
        RECT 50.340 28.510 51.580 28.740 ;
        RECT 53.515 28.740 53.775 29.620 ;
        RECT 54.015 28.900 54.245 29.790 ;
        RECT 54.805 28.900 55.035 29.790 ;
        RECT 55.395 28.900 55.625 29.790 ;
        RECT 56.185 28.900 56.415 29.865 ;
        RECT 59.325 29.790 59.585 30.110 ;
        RECT 60.115 29.790 60.375 30.110 ;
        RECT 60.705 29.790 60.965 30.110 ;
        RECT 61.510 30.035 61.740 31.345 ;
        RECT 61.930 30.475 62.190 31.550 ;
        RECT 62.350 30.035 62.520 31.975 ;
        RECT 61.510 29.865 62.520 30.035 ;
        RECT 62.665 29.865 63.020 31.975 ;
        RECT 63.400 32.250 63.755 34.445 ;
        RECT 64.675 34.380 64.905 35.345 ;
        RECT 65.465 34.470 65.695 35.345 ;
        RECT 66.055 34.470 66.285 35.345 ;
        RECT 66.845 34.470 67.075 35.345 ;
        RECT 67.315 34.715 67.575 35.505 ;
        RECT 69.500 35.505 70.740 35.735 ;
        RECT 71.660 35.505 72.900 35.735 ;
        RECT 69.500 34.810 69.760 35.505 ;
        RECT 63.895 34.210 64.905 34.380 ;
        RECT 63.895 32.250 64.065 34.210 ;
        RECT 64.225 32.695 64.485 33.830 ;
        RECT 64.675 32.900 64.905 34.210 ;
        RECT 65.450 34.150 65.710 34.470 ;
        RECT 66.040 34.150 66.300 34.470 ;
        RECT 66.830 34.150 67.090 34.470 ;
        RECT 65.465 32.900 65.695 34.150 ;
        RECT 66.055 32.900 66.285 34.150 ;
        RECT 66.845 32.900 67.075 34.150 ;
        RECT 67.315 32.695 67.575 33.200 ;
        RECT 64.225 32.465 65.415 32.695 ;
        RECT 66.335 32.465 67.575 32.695 ;
        RECT 68.000 32.250 68.355 34.440 ;
        RECT 63.400 31.975 64.065 32.250 ;
        RECT 67.685 31.975 68.355 32.250 ;
        RECT 63.400 29.870 63.755 31.975 ;
        RECT 64.175 31.550 65.415 31.780 ;
        RECT 66.335 31.550 67.525 31.780 ;
        RECT 64.175 31.125 64.435 31.550 ;
        RECT 64.675 30.110 64.905 31.345 ;
        RECT 65.465 30.110 65.695 31.345 ;
        RECT 66.055 30.110 66.285 31.345 ;
        RECT 56.655 28.740 56.915 29.530 ;
        RECT 53.515 28.510 54.755 28.740 ;
        RECT 55.675 28.510 56.915 28.740 ;
        RECT 58.840 28.740 59.100 29.620 ;
        RECT 59.340 28.900 59.570 29.790 ;
        RECT 60.130 28.900 60.360 29.790 ;
        RECT 60.720 28.900 60.950 29.790 ;
        RECT 61.510 28.900 61.740 29.865 ;
        RECT 64.660 29.790 64.920 30.110 ;
        RECT 65.450 29.790 65.710 30.110 ;
        RECT 66.040 29.790 66.300 30.110 ;
        RECT 66.845 30.035 67.075 31.345 ;
        RECT 67.265 30.475 67.525 31.550 ;
        RECT 67.685 30.035 67.855 31.975 ;
        RECT 66.845 29.865 67.855 30.035 ;
        RECT 68.000 29.865 68.355 31.975 ;
        RECT 68.725 32.250 69.080 34.445 ;
        RECT 70.000 34.380 70.230 35.345 ;
        RECT 70.790 34.470 71.020 35.345 ;
        RECT 71.380 34.470 71.610 35.345 ;
        RECT 72.170 34.470 72.400 35.345 ;
        RECT 72.640 34.715 72.900 35.505 ;
        RECT 74.835 35.505 76.075 35.735 ;
        RECT 76.995 35.505 78.235 35.735 ;
        RECT 74.835 34.810 75.095 35.505 ;
        RECT 69.220 34.210 70.230 34.380 ;
        RECT 69.220 32.250 69.390 34.210 ;
        RECT 69.550 32.695 69.810 33.830 ;
        RECT 70.000 32.900 70.230 34.210 ;
        RECT 70.775 34.150 71.035 34.470 ;
        RECT 71.365 34.150 71.625 34.470 ;
        RECT 72.155 34.150 72.415 34.470 ;
        RECT 70.790 32.900 71.020 34.150 ;
        RECT 71.380 32.900 71.610 34.150 ;
        RECT 72.170 32.900 72.400 34.150 ;
        RECT 72.640 32.695 72.900 33.200 ;
        RECT 69.550 32.465 70.740 32.695 ;
        RECT 71.660 32.465 72.900 32.695 ;
        RECT 73.325 32.250 73.680 34.440 ;
        RECT 68.725 31.975 69.390 32.250 ;
        RECT 73.010 31.975 73.680 32.250 ;
        RECT 68.725 29.870 69.080 31.975 ;
        RECT 69.500 31.550 70.740 31.780 ;
        RECT 71.660 31.550 72.850 31.780 ;
        RECT 69.500 31.125 69.760 31.550 ;
        RECT 70.000 30.110 70.230 31.345 ;
        RECT 70.790 30.110 71.020 31.345 ;
        RECT 71.380 30.110 71.610 31.345 ;
        RECT 61.980 28.740 62.240 29.530 ;
        RECT 58.840 28.510 60.080 28.740 ;
        RECT 61.000 28.510 62.240 28.740 ;
        RECT 64.175 28.740 64.435 29.620 ;
        RECT 64.675 28.900 64.905 29.790 ;
        RECT 65.465 28.900 65.695 29.790 ;
        RECT 66.055 28.900 66.285 29.790 ;
        RECT 66.845 28.900 67.075 29.865 ;
        RECT 69.985 29.790 70.245 30.110 ;
        RECT 70.775 29.790 71.035 30.110 ;
        RECT 71.365 29.790 71.625 30.110 ;
        RECT 72.170 30.035 72.400 31.345 ;
        RECT 72.590 30.475 72.850 31.550 ;
        RECT 73.010 30.035 73.180 31.975 ;
        RECT 72.170 29.865 73.180 30.035 ;
        RECT 73.325 29.865 73.680 31.975 ;
        RECT 74.060 32.250 74.415 34.445 ;
        RECT 75.335 34.380 75.565 35.345 ;
        RECT 76.125 34.470 76.355 35.345 ;
        RECT 76.715 34.470 76.945 35.345 ;
        RECT 77.505 34.470 77.735 35.345 ;
        RECT 77.975 34.715 78.235 35.505 ;
        RECT 80.160 35.505 81.400 35.735 ;
        RECT 82.320 35.505 83.560 35.735 ;
        RECT 80.160 34.810 80.420 35.505 ;
        RECT 74.555 34.210 75.565 34.380 ;
        RECT 74.555 32.250 74.725 34.210 ;
        RECT 74.885 32.695 75.145 33.830 ;
        RECT 75.335 32.900 75.565 34.210 ;
        RECT 76.110 34.150 76.370 34.470 ;
        RECT 76.700 34.150 76.960 34.470 ;
        RECT 77.490 34.150 77.750 34.470 ;
        RECT 76.125 32.900 76.355 34.150 ;
        RECT 76.715 32.900 76.945 34.150 ;
        RECT 77.505 32.900 77.735 34.150 ;
        RECT 77.975 32.695 78.235 33.200 ;
        RECT 74.885 32.465 76.075 32.695 ;
        RECT 76.995 32.465 78.235 32.695 ;
        RECT 78.660 32.250 79.015 34.440 ;
        RECT 74.060 31.975 74.725 32.250 ;
        RECT 78.345 31.975 79.015 32.250 ;
        RECT 74.060 29.870 74.415 31.975 ;
        RECT 74.835 31.550 76.075 31.780 ;
        RECT 76.995 31.550 78.185 31.780 ;
        RECT 74.835 31.125 75.095 31.550 ;
        RECT 75.335 30.110 75.565 31.345 ;
        RECT 76.125 30.110 76.355 31.345 ;
        RECT 76.715 30.110 76.945 31.345 ;
        RECT 67.315 28.740 67.575 29.530 ;
        RECT 64.175 28.510 65.415 28.740 ;
        RECT 66.335 28.510 67.575 28.740 ;
        RECT 69.500 28.740 69.760 29.620 ;
        RECT 70.000 28.900 70.230 29.790 ;
        RECT 70.790 28.900 71.020 29.790 ;
        RECT 71.380 28.900 71.610 29.790 ;
        RECT 72.170 28.900 72.400 29.865 ;
        RECT 75.320 29.790 75.580 30.110 ;
        RECT 76.110 29.790 76.370 30.110 ;
        RECT 76.700 29.790 76.960 30.110 ;
        RECT 77.505 30.035 77.735 31.345 ;
        RECT 77.925 30.475 78.185 31.550 ;
        RECT 78.345 30.035 78.515 31.975 ;
        RECT 77.505 29.865 78.515 30.035 ;
        RECT 78.660 29.865 79.015 31.975 ;
        RECT 79.385 32.250 79.740 34.445 ;
        RECT 80.660 34.380 80.890 35.345 ;
        RECT 81.450 34.470 81.680 35.345 ;
        RECT 82.040 34.470 82.270 35.345 ;
        RECT 82.830 34.470 83.060 35.345 ;
        RECT 83.300 34.715 83.560 35.505 ;
        RECT 85.495 35.505 86.735 35.735 ;
        RECT 87.655 35.505 88.895 35.735 ;
        RECT 85.495 34.810 85.755 35.505 ;
        RECT 79.880 34.210 80.890 34.380 ;
        RECT 79.880 32.250 80.050 34.210 ;
        RECT 80.210 32.695 80.470 33.830 ;
        RECT 80.660 32.900 80.890 34.210 ;
        RECT 81.435 34.150 81.695 34.470 ;
        RECT 82.025 34.150 82.285 34.470 ;
        RECT 82.815 34.150 83.075 34.470 ;
        RECT 81.450 32.900 81.680 34.150 ;
        RECT 82.040 32.900 82.270 34.150 ;
        RECT 82.830 32.900 83.060 34.150 ;
        RECT 83.300 32.695 83.560 33.200 ;
        RECT 80.210 32.465 81.400 32.695 ;
        RECT 82.320 32.465 83.560 32.695 ;
        RECT 83.985 32.250 84.340 34.440 ;
        RECT 79.385 31.975 80.050 32.250 ;
        RECT 83.670 31.975 84.340 32.250 ;
        RECT 79.385 29.870 79.740 31.975 ;
        RECT 80.160 31.550 81.400 31.780 ;
        RECT 82.320 31.550 83.510 31.780 ;
        RECT 80.160 31.125 80.420 31.550 ;
        RECT 80.660 30.110 80.890 31.345 ;
        RECT 81.450 30.110 81.680 31.345 ;
        RECT 82.040 30.110 82.270 31.345 ;
        RECT 72.640 28.740 72.900 29.530 ;
        RECT 69.500 28.510 70.740 28.740 ;
        RECT 71.660 28.510 72.900 28.740 ;
        RECT 74.835 28.740 75.095 29.620 ;
        RECT 75.335 28.900 75.565 29.790 ;
        RECT 76.125 28.900 76.355 29.790 ;
        RECT 76.715 28.900 76.945 29.790 ;
        RECT 77.505 28.900 77.735 29.865 ;
        RECT 80.645 29.790 80.905 30.110 ;
        RECT 81.435 29.790 81.695 30.110 ;
        RECT 82.025 29.790 82.285 30.110 ;
        RECT 82.830 30.035 83.060 31.345 ;
        RECT 83.250 30.475 83.510 31.550 ;
        RECT 83.670 30.035 83.840 31.975 ;
        RECT 82.830 29.865 83.840 30.035 ;
        RECT 83.985 29.865 84.340 31.975 ;
        RECT 84.720 32.250 85.075 34.445 ;
        RECT 85.995 34.380 86.225 35.345 ;
        RECT 86.785 34.470 87.015 35.345 ;
        RECT 87.375 34.470 87.605 35.345 ;
        RECT 88.165 34.470 88.395 35.345 ;
        RECT 88.635 34.715 88.895 35.505 ;
        RECT 90.820 35.505 92.060 35.735 ;
        RECT 92.980 35.505 94.220 35.735 ;
        RECT 90.820 34.810 91.080 35.505 ;
        RECT 85.215 34.210 86.225 34.380 ;
        RECT 85.215 32.250 85.385 34.210 ;
        RECT 85.545 32.695 85.805 33.830 ;
        RECT 85.995 32.900 86.225 34.210 ;
        RECT 86.770 34.150 87.030 34.470 ;
        RECT 87.360 34.150 87.620 34.470 ;
        RECT 88.150 34.150 88.410 34.470 ;
        RECT 86.785 32.900 87.015 34.150 ;
        RECT 87.375 32.900 87.605 34.150 ;
        RECT 88.165 32.900 88.395 34.150 ;
        RECT 88.635 32.695 88.895 33.200 ;
        RECT 85.545 32.465 86.735 32.695 ;
        RECT 87.655 32.465 88.895 32.695 ;
        RECT 89.320 32.250 89.675 34.440 ;
        RECT 84.720 31.975 85.385 32.250 ;
        RECT 89.005 31.975 89.675 32.250 ;
        RECT 84.720 29.870 85.075 31.975 ;
        RECT 85.495 31.550 86.735 31.780 ;
        RECT 87.655 31.550 88.845 31.780 ;
        RECT 85.495 31.125 85.755 31.550 ;
        RECT 85.995 30.110 86.225 31.345 ;
        RECT 86.785 30.110 87.015 31.345 ;
        RECT 87.375 30.110 87.605 31.345 ;
        RECT 77.975 28.740 78.235 29.530 ;
        RECT 74.835 28.510 76.075 28.740 ;
        RECT 76.995 28.510 78.235 28.740 ;
        RECT 80.160 28.740 80.420 29.620 ;
        RECT 80.660 28.900 80.890 29.790 ;
        RECT 81.450 28.900 81.680 29.790 ;
        RECT 82.040 28.900 82.270 29.790 ;
        RECT 82.830 28.900 83.060 29.865 ;
        RECT 85.980 29.790 86.240 30.110 ;
        RECT 86.770 29.790 87.030 30.110 ;
        RECT 87.360 29.790 87.620 30.110 ;
        RECT 88.165 30.035 88.395 31.345 ;
        RECT 88.585 30.475 88.845 31.550 ;
        RECT 89.005 30.035 89.175 31.975 ;
        RECT 88.165 29.865 89.175 30.035 ;
        RECT 89.320 29.865 89.675 31.975 ;
        RECT 90.045 32.250 90.400 34.445 ;
        RECT 91.320 34.380 91.550 35.345 ;
        RECT 92.110 34.470 92.340 35.345 ;
        RECT 92.700 34.470 92.930 35.345 ;
        RECT 93.490 34.470 93.720 35.345 ;
        RECT 93.960 34.715 94.220 35.505 ;
        RECT 96.155 35.505 97.395 35.735 ;
        RECT 98.315 35.505 99.555 35.735 ;
        RECT 96.155 34.810 96.415 35.505 ;
        RECT 90.540 34.210 91.550 34.380 ;
        RECT 90.540 32.250 90.710 34.210 ;
        RECT 90.870 32.695 91.130 33.830 ;
        RECT 91.320 32.900 91.550 34.210 ;
        RECT 92.095 34.150 92.355 34.470 ;
        RECT 92.685 34.150 92.945 34.470 ;
        RECT 93.475 34.150 93.735 34.470 ;
        RECT 92.110 32.900 92.340 34.150 ;
        RECT 92.700 32.900 92.930 34.150 ;
        RECT 93.490 32.900 93.720 34.150 ;
        RECT 93.960 32.695 94.220 33.200 ;
        RECT 90.870 32.465 92.060 32.695 ;
        RECT 92.980 32.465 94.220 32.695 ;
        RECT 94.645 32.250 95.000 34.440 ;
        RECT 90.045 31.975 90.710 32.250 ;
        RECT 94.330 31.975 95.000 32.250 ;
        RECT 90.045 29.870 90.400 31.975 ;
        RECT 90.820 31.550 92.060 31.780 ;
        RECT 92.980 31.550 94.170 31.780 ;
        RECT 90.820 31.125 91.080 31.550 ;
        RECT 91.320 30.110 91.550 31.345 ;
        RECT 92.110 30.110 92.340 31.345 ;
        RECT 92.700 30.110 92.930 31.345 ;
        RECT 83.300 28.740 83.560 29.530 ;
        RECT 80.160 28.510 81.400 28.740 ;
        RECT 82.320 28.510 83.560 28.740 ;
        RECT 85.495 28.740 85.755 29.620 ;
        RECT 85.995 28.900 86.225 29.790 ;
        RECT 86.785 28.900 87.015 29.790 ;
        RECT 87.375 28.900 87.605 29.790 ;
        RECT 88.165 28.900 88.395 29.865 ;
        RECT 91.305 29.790 91.565 30.110 ;
        RECT 92.095 29.790 92.355 30.110 ;
        RECT 92.685 29.790 92.945 30.110 ;
        RECT 93.490 30.035 93.720 31.345 ;
        RECT 93.910 30.475 94.170 31.550 ;
        RECT 94.330 30.035 94.500 31.975 ;
        RECT 93.490 29.865 94.500 30.035 ;
        RECT 94.645 29.865 95.000 31.975 ;
        RECT 95.380 32.250 95.735 34.445 ;
        RECT 96.655 34.380 96.885 35.345 ;
        RECT 97.445 34.470 97.675 35.345 ;
        RECT 98.035 34.470 98.265 35.345 ;
        RECT 98.825 34.470 99.055 35.345 ;
        RECT 99.295 34.715 99.555 35.505 ;
        RECT 101.480 35.505 102.720 35.735 ;
        RECT 103.640 35.505 104.880 35.735 ;
        RECT 101.480 34.810 101.740 35.505 ;
        RECT 95.875 34.210 96.885 34.380 ;
        RECT 95.875 32.250 96.045 34.210 ;
        RECT 96.205 32.695 96.465 33.830 ;
        RECT 96.655 32.900 96.885 34.210 ;
        RECT 97.430 34.150 97.690 34.470 ;
        RECT 98.020 34.150 98.280 34.470 ;
        RECT 98.810 34.150 99.070 34.470 ;
        RECT 97.445 32.900 97.675 34.150 ;
        RECT 98.035 32.900 98.265 34.150 ;
        RECT 98.825 32.900 99.055 34.150 ;
        RECT 99.295 32.695 99.555 33.200 ;
        RECT 96.205 32.465 97.395 32.695 ;
        RECT 98.315 32.465 99.555 32.695 ;
        RECT 99.980 32.250 100.335 34.440 ;
        RECT 95.380 31.975 96.045 32.250 ;
        RECT 99.665 31.975 100.335 32.250 ;
        RECT 95.380 29.870 95.735 31.975 ;
        RECT 96.155 31.550 97.395 31.780 ;
        RECT 98.315 31.550 99.505 31.780 ;
        RECT 96.155 31.125 96.415 31.550 ;
        RECT 96.655 30.110 96.885 31.345 ;
        RECT 97.445 30.110 97.675 31.345 ;
        RECT 98.035 30.110 98.265 31.345 ;
        RECT 88.635 28.740 88.895 29.530 ;
        RECT 85.495 28.510 86.735 28.740 ;
        RECT 87.655 28.510 88.895 28.740 ;
        RECT 90.820 28.740 91.080 29.620 ;
        RECT 91.320 28.900 91.550 29.790 ;
        RECT 92.110 28.900 92.340 29.790 ;
        RECT 92.700 28.900 92.930 29.790 ;
        RECT 93.490 28.900 93.720 29.865 ;
        RECT 96.640 29.790 96.900 30.110 ;
        RECT 97.430 29.790 97.690 30.110 ;
        RECT 98.020 29.790 98.280 30.110 ;
        RECT 98.825 30.035 99.055 31.345 ;
        RECT 99.245 30.475 99.505 31.550 ;
        RECT 99.665 30.035 99.835 31.975 ;
        RECT 98.825 29.865 99.835 30.035 ;
        RECT 99.980 29.865 100.335 31.975 ;
        RECT 100.705 32.250 101.060 34.445 ;
        RECT 101.980 34.380 102.210 35.345 ;
        RECT 102.770 34.470 103.000 35.345 ;
        RECT 103.360 34.470 103.590 35.345 ;
        RECT 104.150 34.470 104.380 35.345 ;
        RECT 104.620 34.715 104.880 35.505 ;
        RECT 106.815 35.505 108.055 35.735 ;
        RECT 108.975 35.505 110.215 35.735 ;
        RECT 106.815 34.810 107.075 35.505 ;
        RECT 101.200 34.210 102.210 34.380 ;
        RECT 101.200 32.250 101.370 34.210 ;
        RECT 101.530 32.695 101.790 33.830 ;
        RECT 101.980 32.900 102.210 34.210 ;
        RECT 102.755 34.150 103.015 34.470 ;
        RECT 103.345 34.150 103.605 34.470 ;
        RECT 104.135 34.150 104.395 34.470 ;
        RECT 102.770 32.900 103.000 34.150 ;
        RECT 103.360 32.900 103.590 34.150 ;
        RECT 104.150 32.900 104.380 34.150 ;
        RECT 104.620 32.695 104.880 33.200 ;
        RECT 101.530 32.465 102.720 32.695 ;
        RECT 103.640 32.465 104.880 32.695 ;
        RECT 105.305 32.250 105.660 34.440 ;
        RECT 100.705 31.975 101.370 32.250 ;
        RECT 104.990 31.975 105.660 32.250 ;
        RECT 100.705 29.870 101.060 31.975 ;
        RECT 101.480 31.550 102.720 31.780 ;
        RECT 103.640 31.550 104.830 31.780 ;
        RECT 101.480 31.125 101.740 31.550 ;
        RECT 101.980 30.110 102.210 31.345 ;
        RECT 102.770 30.110 103.000 31.345 ;
        RECT 103.360 30.110 103.590 31.345 ;
        RECT 93.960 28.740 94.220 29.530 ;
        RECT 90.820 28.510 92.060 28.740 ;
        RECT 92.980 28.510 94.220 28.740 ;
        RECT 96.155 28.740 96.415 29.620 ;
        RECT 96.655 28.900 96.885 29.790 ;
        RECT 97.445 28.900 97.675 29.790 ;
        RECT 98.035 28.900 98.265 29.790 ;
        RECT 98.825 28.900 99.055 29.865 ;
        RECT 101.965 29.790 102.225 30.110 ;
        RECT 102.755 29.790 103.015 30.110 ;
        RECT 103.345 29.790 103.605 30.110 ;
        RECT 104.150 30.035 104.380 31.345 ;
        RECT 104.570 30.475 104.830 31.550 ;
        RECT 104.990 30.035 105.160 31.975 ;
        RECT 104.150 29.865 105.160 30.035 ;
        RECT 105.305 29.865 105.660 31.975 ;
        RECT 106.040 32.250 106.395 34.445 ;
        RECT 107.315 34.380 107.545 35.345 ;
        RECT 108.105 34.470 108.335 35.345 ;
        RECT 108.695 34.470 108.925 35.345 ;
        RECT 109.485 34.470 109.715 35.345 ;
        RECT 109.955 34.715 110.215 35.505 ;
        RECT 112.140 35.505 113.380 35.735 ;
        RECT 114.300 35.505 115.540 35.735 ;
        RECT 112.140 34.810 112.400 35.505 ;
        RECT 106.535 34.210 107.545 34.380 ;
        RECT 106.535 32.250 106.705 34.210 ;
        RECT 106.865 32.695 107.125 33.830 ;
        RECT 107.315 32.900 107.545 34.210 ;
        RECT 108.090 34.150 108.350 34.470 ;
        RECT 108.680 34.150 108.940 34.470 ;
        RECT 109.470 34.150 109.730 34.470 ;
        RECT 108.105 32.900 108.335 34.150 ;
        RECT 108.695 32.900 108.925 34.150 ;
        RECT 109.485 32.900 109.715 34.150 ;
        RECT 109.955 32.695 110.215 33.200 ;
        RECT 106.865 32.465 108.055 32.695 ;
        RECT 108.975 32.465 110.215 32.695 ;
        RECT 110.640 32.250 110.995 34.440 ;
        RECT 106.040 31.975 106.705 32.250 ;
        RECT 110.325 31.975 110.995 32.250 ;
        RECT 106.040 29.870 106.395 31.975 ;
        RECT 106.815 31.550 108.055 31.780 ;
        RECT 108.975 31.550 110.165 31.780 ;
        RECT 106.815 31.125 107.075 31.550 ;
        RECT 107.315 30.110 107.545 31.345 ;
        RECT 108.105 30.110 108.335 31.345 ;
        RECT 108.695 30.110 108.925 31.345 ;
        RECT 99.295 28.740 99.555 29.530 ;
        RECT 96.155 28.510 97.395 28.740 ;
        RECT 98.315 28.510 99.555 28.740 ;
        RECT 101.480 28.740 101.740 29.620 ;
        RECT 101.980 28.900 102.210 29.790 ;
        RECT 102.770 28.900 103.000 29.790 ;
        RECT 103.360 28.900 103.590 29.790 ;
        RECT 104.150 28.900 104.380 29.865 ;
        RECT 107.300 29.790 107.560 30.110 ;
        RECT 108.090 29.790 108.350 30.110 ;
        RECT 108.680 29.790 108.940 30.110 ;
        RECT 109.485 30.035 109.715 31.345 ;
        RECT 109.905 30.475 110.165 31.550 ;
        RECT 110.325 30.035 110.495 31.975 ;
        RECT 109.485 29.865 110.495 30.035 ;
        RECT 110.640 29.865 110.995 31.975 ;
        RECT 111.365 32.250 111.720 34.445 ;
        RECT 112.640 34.380 112.870 35.345 ;
        RECT 113.430 34.470 113.660 35.345 ;
        RECT 114.020 34.470 114.250 35.345 ;
        RECT 114.810 34.470 115.040 35.345 ;
        RECT 115.280 34.715 115.540 35.505 ;
        RECT 117.475 35.505 118.715 35.735 ;
        RECT 119.635 35.505 120.875 35.735 ;
        RECT 117.475 34.810 117.735 35.505 ;
        RECT 111.860 34.210 112.870 34.380 ;
        RECT 111.860 32.250 112.030 34.210 ;
        RECT 112.190 32.695 112.450 33.830 ;
        RECT 112.640 32.900 112.870 34.210 ;
        RECT 113.415 34.150 113.675 34.470 ;
        RECT 114.005 34.150 114.265 34.470 ;
        RECT 114.795 34.150 115.055 34.470 ;
        RECT 113.430 32.900 113.660 34.150 ;
        RECT 114.020 32.900 114.250 34.150 ;
        RECT 114.810 32.900 115.040 34.150 ;
        RECT 115.280 32.695 115.540 33.200 ;
        RECT 112.190 32.465 113.380 32.695 ;
        RECT 114.300 32.465 115.540 32.695 ;
        RECT 115.965 32.250 116.320 34.440 ;
        RECT 111.365 31.975 112.030 32.250 ;
        RECT 115.650 31.975 116.320 32.250 ;
        RECT 111.365 29.870 111.720 31.975 ;
        RECT 112.140 31.550 113.380 31.780 ;
        RECT 114.300 31.550 115.490 31.780 ;
        RECT 112.140 31.125 112.400 31.550 ;
        RECT 112.640 30.110 112.870 31.345 ;
        RECT 113.430 30.110 113.660 31.345 ;
        RECT 114.020 30.110 114.250 31.345 ;
        RECT 104.620 28.740 104.880 29.530 ;
        RECT 101.480 28.510 102.720 28.740 ;
        RECT 103.640 28.510 104.880 28.740 ;
        RECT 106.815 28.740 107.075 29.620 ;
        RECT 107.315 28.900 107.545 29.790 ;
        RECT 108.105 28.900 108.335 29.790 ;
        RECT 108.695 28.900 108.925 29.790 ;
        RECT 109.485 28.900 109.715 29.865 ;
        RECT 112.625 29.790 112.885 30.110 ;
        RECT 113.415 29.790 113.675 30.110 ;
        RECT 114.005 29.790 114.265 30.110 ;
        RECT 114.810 30.035 115.040 31.345 ;
        RECT 115.230 30.475 115.490 31.550 ;
        RECT 115.650 30.035 115.820 31.975 ;
        RECT 114.810 29.865 115.820 30.035 ;
        RECT 115.965 29.865 116.320 31.975 ;
        RECT 116.700 32.250 117.055 34.445 ;
        RECT 117.975 34.380 118.205 35.345 ;
        RECT 118.765 34.470 118.995 35.345 ;
        RECT 119.355 34.470 119.585 35.345 ;
        RECT 120.145 34.470 120.375 35.345 ;
        RECT 120.615 34.715 120.875 35.505 ;
        RECT 117.195 34.210 118.205 34.380 ;
        RECT 117.195 32.250 117.365 34.210 ;
        RECT 117.525 32.695 117.785 33.830 ;
        RECT 117.975 32.900 118.205 34.210 ;
        RECT 118.750 34.150 119.010 34.470 ;
        RECT 119.340 34.150 119.600 34.470 ;
        RECT 120.130 34.150 120.390 34.470 ;
        RECT 118.765 32.900 118.995 34.150 ;
        RECT 119.355 32.900 119.585 34.150 ;
        RECT 120.145 32.900 120.375 34.150 ;
        RECT 120.615 32.695 120.875 33.200 ;
        RECT 117.525 32.465 118.715 32.695 ;
        RECT 119.635 32.465 120.875 32.695 ;
        RECT 121.300 32.250 121.655 34.440 ;
        RECT 116.700 31.975 117.365 32.250 ;
        RECT 120.985 31.975 121.655 32.250 ;
        RECT 116.700 29.870 117.055 31.975 ;
        RECT 117.475 31.550 118.715 31.780 ;
        RECT 119.635 31.550 120.825 31.780 ;
        RECT 117.475 31.125 117.735 31.550 ;
        RECT 117.975 30.110 118.205 31.345 ;
        RECT 118.765 30.110 118.995 31.345 ;
        RECT 119.355 30.110 119.585 31.345 ;
        RECT 109.955 28.740 110.215 29.530 ;
        RECT 106.815 28.510 108.055 28.740 ;
        RECT 108.975 28.510 110.215 28.740 ;
        RECT 112.140 28.740 112.400 29.620 ;
        RECT 112.640 28.900 112.870 29.790 ;
        RECT 113.430 28.900 113.660 29.790 ;
        RECT 114.020 28.900 114.250 29.790 ;
        RECT 114.810 28.900 115.040 29.865 ;
        RECT 117.960 29.790 118.220 30.110 ;
        RECT 118.750 29.790 119.010 30.110 ;
        RECT 119.340 29.790 119.600 30.110 ;
        RECT 120.145 30.035 120.375 31.345 ;
        RECT 120.565 30.475 120.825 31.550 ;
        RECT 120.985 30.035 121.155 31.975 ;
        RECT 120.145 29.865 121.155 30.035 ;
        RECT 121.300 29.865 121.655 31.975 ;
        RECT 122.025 32.250 122.380 34.460 ;
        RECT 123.300 34.380 123.530 35.345 ;
        RECT 124.090 34.470 124.320 35.345 ;
        RECT 124.680 34.470 124.910 35.345 ;
        RECT 125.470 34.470 125.700 35.345 ;
        RECT 122.520 34.210 123.530 34.380 ;
        RECT 122.520 32.250 122.690 34.210 ;
        RECT 123.300 32.900 123.530 34.210 ;
        RECT 124.075 34.150 124.335 34.470 ;
        RECT 124.665 34.150 124.925 34.470 ;
        RECT 125.455 34.150 125.715 34.470 ;
        RECT 124.090 32.900 124.320 34.150 ;
        RECT 124.680 32.900 124.910 34.150 ;
        RECT 125.470 32.900 125.700 34.150 ;
        RECT 126.625 32.250 126.980 34.460 ;
        RECT 122.025 31.975 122.690 32.250 ;
        RECT 126.310 31.975 126.980 32.250 ;
        RECT 122.025 29.885 122.380 31.975 ;
        RECT 123.300 30.110 123.530 31.345 ;
        RECT 124.090 30.110 124.320 31.345 ;
        RECT 124.680 30.110 124.910 31.345 ;
        RECT 115.280 28.740 115.540 29.530 ;
        RECT 112.140 28.510 113.380 28.740 ;
        RECT 114.300 28.510 115.540 28.740 ;
        RECT 117.475 28.740 117.735 29.620 ;
        RECT 117.975 28.900 118.205 29.790 ;
        RECT 118.765 28.900 118.995 29.790 ;
        RECT 119.355 28.900 119.585 29.790 ;
        RECT 120.145 28.900 120.375 29.865 ;
        RECT 123.285 29.790 123.545 30.110 ;
        RECT 124.075 29.790 124.335 30.110 ;
        RECT 124.665 29.790 124.925 30.110 ;
        RECT 125.470 30.035 125.700 31.345 ;
        RECT 126.310 30.035 126.480 31.975 ;
        RECT 125.470 29.865 126.480 30.035 ;
        RECT 126.625 29.885 126.980 31.975 ;
        RECT 120.615 28.740 120.875 29.530 ;
        RECT 123.300 28.900 123.530 29.790 ;
        RECT 124.090 28.900 124.320 29.790 ;
        RECT 124.680 28.900 124.910 29.790 ;
        RECT 125.470 28.900 125.700 29.865 ;
        RECT 117.475 28.510 118.715 28.740 ;
        RECT 119.635 28.510 120.875 28.740 ;
        RECT 16.115 28.160 26.090 28.395 ;
        RECT 10.500 27.720 11.960 28.050 ;
        RECT 10.500 27.500 10.820 27.720 ;
        RECT 12.400 26.975 12.720 27.965 ;
        RECT 14.585 27.720 16.005 28.045 ;
        RECT 19.990 27.590 26.090 28.160 ;
        RECT 37.520 27.970 38.760 28.200 ;
        RECT 39.680 27.970 40.920 28.200 ;
        RECT 16.115 27.355 26.090 27.590 ;
        RECT 12.425 26.960 12.715 26.975 ;
        RECT 26.905 24.975 27.165 24.980 ;
        RECT 10.510 23.455 10.810 24.905 ;
        RECT 15.985 24.740 27.225 24.975 ;
        RECT 11.745 24.355 13.345 24.645 ;
        RECT 14.165 24.355 20.945 24.590 ;
        RECT 16.040 24.170 17.645 24.200 ;
        RECT 21.425 24.170 27.225 24.740 ;
        RECT 15.985 23.935 27.225 24.170 ;
        RECT 31.420 24.715 31.775 26.925 ;
        RECT 32.695 26.845 32.925 27.810 ;
        RECT 33.485 26.935 33.715 27.810 ;
        RECT 34.075 26.935 34.305 27.810 ;
        RECT 34.865 26.935 35.095 27.810 ;
        RECT 37.520 27.275 37.780 27.970 ;
        RECT 31.915 26.675 32.925 26.845 ;
        RECT 31.915 24.715 32.085 26.675 ;
        RECT 32.695 25.365 32.925 26.675 ;
        RECT 33.470 26.615 33.730 26.935 ;
        RECT 34.060 26.615 34.320 26.935 ;
        RECT 34.850 26.615 35.110 26.935 ;
        RECT 33.485 25.365 33.715 26.615 ;
        RECT 34.075 25.365 34.305 26.615 ;
        RECT 34.865 25.365 35.095 26.615 ;
        RECT 36.020 24.715 36.375 26.925 ;
        RECT 31.420 24.440 32.085 24.715 ;
        RECT 35.705 24.440 36.375 24.715 ;
        RECT 16.040 23.910 17.645 23.935 ;
        RECT 31.420 22.350 31.775 24.440 ;
        RECT 32.695 22.575 32.925 23.810 ;
        RECT 33.485 22.575 33.715 23.810 ;
        RECT 34.075 22.575 34.305 23.810 ;
        RECT 32.680 22.255 32.940 22.575 ;
        RECT 33.470 22.255 33.730 22.575 ;
        RECT 34.060 22.255 34.320 22.575 ;
        RECT 34.865 22.500 35.095 23.810 ;
        RECT 35.705 22.500 35.875 24.440 ;
        RECT 34.865 22.330 35.875 22.500 ;
        RECT 36.020 22.350 36.375 24.440 ;
        RECT 36.745 24.715 37.100 26.910 ;
        RECT 38.020 26.845 38.250 27.810 ;
        RECT 38.810 26.935 39.040 27.810 ;
        RECT 39.400 26.935 39.630 27.810 ;
        RECT 40.190 26.935 40.420 27.810 ;
        RECT 40.660 27.180 40.920 27.970 ;
        RECT 42.855 27.970 44.095 28.200 ;
        RECT 45.015 27.970 46.255 28.200 ;
        RECT 42.855 27.275 43.115 27.970 ;
        RECT 37.240 26.675 38.250 26.845 ;
        RECT 37.240 24.715 37.410 26.675 ;
        RECT 37.570 25.160 37.830 26.295 ;
        RECT 38.020 25.365 38.250 26.675 ;
        RECT 38.795 26.615 39.055 26.935 ;
        RECT 39.385 26.615 39.645 26.935 ;
        RECT 40.175 26.615 40.435 26.935 ;
        RECT 38.810 25.365 39.040 26.615 ;
        RECT 39.400 25.365 39.630 26.615 ;
        RECT 40.190 25.365 40.420 26.615 ;
        RECT 40.660 25.160 40.920 25.665 ;
        RECT 37.570 24.930 38.760 25.160 ;
        RECT 39.680 24.930 40.920 25.160 ;
        RECT 41.345 24.715 41.700 26.905 ;
        RECT 36.745 24.440 37.410 24.715 ;
        RECT 41.030 24.440 41.700 24.715 ;
        RECT 36.745 22.335 37.100 24.440 ;
        RECT 37.520 24.015 38.760 24.245 ;
        RECT 39.680 24.015 40.870 24.245 ;
        RECT 37.520 23.590 37.780 24.015 ;
        RECT 38.020 22.575 38.250 23.810 ;
        RECT 38.810 22.575 39.040 23.810 ;
        RECT 39.400 22.575 39.630 23.810 ;
        RECT 32.695 21.365 32.925 22.255 ;
        RECT 33.485 21.365 33.715 22.255 ;
        RECT 34.075 21.365 34.305 22.255 ;
        RECT 34.865 21.365 35.095 22.330 ;
        RECT 38.005 22.255 38.265 22.575 ;
        RECT 38.795 22.255 39.055 22.575 ;
        RECT 39.385 22.255 39.645 22.575 ;
        RECT 40.190 22.500 40.420 23.810 ;
        RECT 40.610 22.940 40.870 24.015 ;
        RECT 41.030 22.500 41.200 24.440 ;
        RECT 40.190 22.330 41.200 22.500 ;
        RECT 41.345 22.330 41.700 24.440 ;
        RECT 42.080 24.715 42.435 26.910 ;
        RECT 43.355 26.845 43.585 27.810 ;
        RECT 44.145 26.935 44.375 27.810 ;
        RECT 44.735 26.935 44.965 27.810 ;
        RECT 45.525 26.935 45.755 27.810 ;
        RECT 45.995 27.180 46.255 27.970 ;
        RECT 48.180 27.970 49.420 28.200 ;
        RECT 50.340 27.970 51.580 28.200 ;
        RECT 48.180 27.275 48.440 27.970 ;
        RECT 42.575 26.675 43.585 26.845 ;
        RECT 42.575 24.715 42.745 26.675 ;
        RECT 42.905 25.160 43.165 26.295 ;
        RECT 43.355 25.365 43.585 26.675 ;
        RECT 44.130 26.615 44.390 26.935 ;
        RECT 44.720 26.615 44.980 26.935 ;
        RECT 45.510 26.615 45.770 26.935 ;
        RECT 44.145 25.365 44.375 26.615 ;
        RECT 44.735 25.365 44.965 26.615 ;
        RECT 45.525 25.365 45.755 26.615 ;
        RECT 45.995 25.160 46.255 25.665 ;
        RECT 42.905 24.930 44.095 25.160 ;
        RECT 45.015 24.930 46.255 25.160 ;
        RECT 46.680 24.715 47.035 26.905 ;
        RECT 42.080 24.440 42.745 24.715 ;
        RECT 46.365 24.440 47.035 24.715 ;
        RECT 42.080 22.335 42.435 24.440 ;
        RECT 42.855 24.015 44.095 24.245 ;
        RECT 45.015 24.015 46.205 24.245 ;
        RECT 42.855 23.590 43.115 24.015 ;
        RECT 43.355 22.575 43.585 23.810 ;
        RECT 44.145 22.575 44.375 23.810 ;
        RECT 44.735 22.575 44.965 23.810 ;
        RECT 37.520 21.205 37.780 22.085 ;
        RECT 38.020 21.365 38.250 22.255 ;
        RECT 38.810 21.365 39.040 22.255 ;
        RECT 39.400 21.365 39.630 22.255 ;
        RECT 40.190 21.365 40.420 22.330 ;
        RECT 43.340 22.255 43.600 22.575 ;
        RECT 44.130 22.255 44.390 22.575 ;
        RECT 44.720 22.255 44.980 22.575 ;
        RECT 45.525 22.500 45.755 23.810 ;
        RECT 45.945 22.940 46.205 24.015 ;
        RECT 46.365 22.500 46.535 24.440 ;
        RECT 45.525 22.330 46.535 22.500 ;
        RECT 46.680 22.330 47.035 24.440 ;
        RECT 47.405 24.715 47.760 26.910 ;
        RECT 48.680 26.845 48.910 27.810 ;
        RECT 49.470 26.935 49.700 27.810 ;
        RECT 50.060 26.935 50.290 27.810 ;
        RECT 50.850 26.935 51.080 27.810 ;
        RECT 51.320 27.180 51.580 27.970 ;
        RECT 53.515 27.970 54.755 28.200 ;
        RECT 55.675 27.970 56.915 28.200 ;
        RECT 53.515 27.275 53.775 27.970 ;
        RECT 47.900 26.675 48.910 26.845 ;
        RECT 47.900 24.715 48.070 26.675 ;
        RECT 48.230 25.160 48.490 26.295 ;
        RECT 48.680 25.365 48.910 26.675 ;
        RECT 49.455 26.615 49.715 26.935 ;
        RECT 50.045 26.615 50.305 26.935 ;
        RECT 50.835 26.615 51.095 26.935 ;
        RECT 49.470 25.365 49.700 26.615 ;
        RECT 50.060 25.365 50.290 26.615 ;
        RECT 50.850 25.365 51.080 26.615 ;
        RECT 51.320 25.160 51.580 25.665 ;
        RECT 48.230 24.930 49.420 25.160 ;
        RECT 50.340 24.930 51.580 25.160 ;
        RECT 52.005 24.715 52.360 26.905 ;
        RECT 47.405 24.440 48.070 24.715 ;
        RECT 51.690 24.440 52.360 24.715 ;
        RECT 47.405 22.335 47.760 24.440 ;
        RECT 48.180 24.015 49.420 24.245 ;
        RECT 50.340 24.015 51.530 24.245 ;
        RECT 48.180 23.590 48.440 24.015 ;
        RECT 48.680 22.575 48.910 23.810 ;
        RECT 49.470 22.575 49.700 23.810 ;
        RECT 50.060 22.575 50.290 23.810 ;
        RECT 40.660 21.205 40.920 21.995 ;
        RECT 37.520 20.975 38.760 21.205 ;
        RECT 39.680 20.975 40.920 21.205 ;
        RECT 42.855 21.205 43.115 22.085 ;
        RECT 43.355 21.365 43.585 22.255 ;
        RECT 44.145 21.365 44.375 22.255 ;
        RECT 44.735 21.365 44.965 22.255 ;
        RECT 45.525 21.365 45.755 22.330 ;
        RECT 48.665 22.255 48.925 22.575 ;
        RECT 49.455 22.255 49.715 22.575 ;
        RECT 50.045 22.255 50.305 22.575 ;
        RECT 50.850 22.500 51.080 23.810 ;
        RECT 51.270 22.940 51.530 24.015 ;
        RECT 51.690 22.500 51.860 24.440 ;
        RECT 50.850 22.330 51.860 22.500 ;
        RECT 52.005 22.330 52.360 24.440 ;
        RECT 52.740 24.715 53.095 26.910 ;
        RECT 54.015 26.845 54.245 27.810 ;
        RECT 54.805 26.935 55.035 27.810 ;
        RECT 55.395 26.935 55.625 27.810 ;
        RECT 56.185 26.935 56.415 27.810 ;
        RECT 56.655 27.180 56.915 27.970 ;
        RECT 58.840 27.970 60.080 28.200 ;
        RECT 61.000 27.970 62.240 28.200 ;
        RECT 58.840 27.275 59.100 27.970 ;
        RECT 53.235 26.675 54.245 26.845 ;
        RECT 53.235 24.715 53.405 26.675 ;
        RECT 53.565 25.160 53.825 26.295 ;
        RECT 54.015 25.365 54.245 26.675 ;
        RECT 54.790 26.615 55.050 26.935 ;
        RECT 55.380 26.615 55.640 26.935 ;
        RECT 56.170 26.615 56.430 26.935 ;
        RECT 54.805 25.365 55.035 26.615 ;
        RECT 55.395 25.365 55.625 26.615 ;
        RECT 56.185 25.365 56.415 26.615 ;
        RECT 56.655 25.160 56.915 25.665 ;
        RECT 53.565 24.930 54.755 25.160 ;
        RECT 55.675 24.930 56.915 25.160 ;
        RECT 57.340 24.715 57.695 26.905 ;
        RECT 52.740 24.440 53.405 24.715 ;
        RECT 57.025 24.440 57.695 24.715 ;
        RECT 52.740 22.335 53.095 24.440 ;
        RECT 53.515 24.015 54.755 24.245 ;
        RECT 55.675 24.015 56.865 24.245 ;
        RECT 53.515 23.590 53.775 24.015 ;
        RECT 54.015 22.575 54.245 23.810 ;
        RECT 54.805 22.575 55.035 23.810 ;
        RECT 55.395 22.575 55.625 23.810 ;
        RECT 45.995 21.205 46.255 21.995 ;
        RECT 42.855 20.975 44.095 21.205 ;
        RECT 45.015 20.975 46.255 21.205 ;
        RECT 48.180 21.205 48.440 22.085 ;
        RECT 48.680 21.365 48.910 22.255 ;
        RECT 49.470 21.365 49.700 22.255 ;
        RECT 50.060 21.365 50.290 22.255 ;
        RECT 50.850 21.365 51.080 22.330 ;
        RECT 54.000 22.255 54.260 22.575 ;
        RECT 54.790 22.255 55.050 22.575 ;
        RECT 55.380 22.255 55.640 22.575 ;
        RECT 56.185 22.500 56.415 23.810 ;
        RECT 56.605 22.940 56.865 24.015 ;
        RECT 57.025 22.500 57.195 24.440 ;
        RECT 56.185 22.330 57.195 22.500 ;
        RECT 57.340 22.330 57.695 24.440 ;
        RECT 58.065 24.715 58.420 26.910 ;
        RECT 59.340 26.845 59.570 27.810 ;
        RECT 60.130 26.935 60.360 27.810 ;
        RECT 60.720 26.935 60.950 27.810 ;
        RECT 61.510 26.935 61.740 27.810 ;
        RECT 61.980 27.180 62.240 27.970 ;
        RECT 64.175 27.970 65.415 28.200 ;
        RECT 66.335 27.970 67.575 28.200 ;
        RECT 64.175 27.275 64.435 27.970 ;
        RECT 58.560 26.675 59.570 26.845 ;
        RECT 58.560 24.715 58.730 26.675 ;
        RECT 58.890 25.160 59.150 26.295 ;
        RECT 59.340 25.365 59.570 26.675 ;
        RECT 60.115 26.615 60.375 26.935 ;
        RECT 60.705 26.615 60.965 26.935 ;
        RECT 61.495 26.615 61.755 26.935 ;
        RECT 60.130 25.365 60.360 26.615 ;
        RECT 60.720 25.365 60.950 26.615 ;
        RECT 61.510 25.365 61.740 26.615 ;
        RECT 61.980 25.160 62.240 25.665 ;
        RECT 58.890 24.930 60.080 25.160 ;
        RECT 61.000 24.930 62.240 25.160 ;
        RECT 62.665 24.715 63.020 26.905 ;
        RECT 58.065 24.440 58.730 24.715 ;
        RECT 62.350 24.440 63.020 24.715 ;
        RECT 58.065 22.335 58.420 24.440 ;
        RECT 58.840 24.015 60.080 24.245 ;
        RECT 61.000 24.015 62.190 24.245 ;
        RECT 58.840 23.590 59.100 24.015 ;
        RECT 59.340 22.575 59.570 23.810 ;
        RECT 60.130 22.575 60.360 23.810 ;
        RECT 60.720 22.575 60.950 23.810 ;
        RECT 51.320 21.205 51.580 21.995 ;
        RECT 48.180 20.975 49.420 21.205 ;
        RECT 50.340 20.975 51.580 21.205 ;
        RECT 53.515 21.205 53.775 22.085 ;
        RECT 54.015 21.365 54.245 22.255 ;
        RECT 54.805 21.365 55.035 22.255 ;
        RECT 55.395 21.365 55.625 22.255 ;
        RECT 56.185 21.365 56.415 22.330 ;
        RECT 59.325 22.255 59.585 22.575 ;
        RECT 60.115 22.255 60.375 22.575 ;
        RECT 60.705 22.255 60.965 22.575 ;
        RECT 61.510 22.500 61.740 23.810 ;
        RECT 61.930 22.940 62.190 24.015 ;
        RECT 62.350 22.500 62.520 24.440 ;
        RECT 61.510 22.330 62.520 22.500 ;
        RECT 62.665 22.330 63.020 24.440 ;
        RECT 63.400 24.715 63.755 26.910 ;
        RECT 64.675 26.845 64.905 27.810 ;
        RECT 65.465 26.935 65.695 27.810 ;
        RECT 66.055 26.935 66.285 27.810 ;
        RECT 66.845 26.935 67.075 27.810 ;
        RECT 67.315 27.180 67.575 27.970 ;
        RECT 69.500 27.970 70.740 28.200 ;
        RECT 71.660 27.970 72.900 28.200 ;
        RECT 69.500 27.275 69.760 27.970 ;
        RECT 63.895 26.675 64.905 26.845 ;
        RECT 63.895 24.715 64.065 26.675 ;
        RECT 64.225 25.160 64.485 26.295 ;
        RECT 64.675 25.365 64.905 26.675 ;
        RECT 65.450 26.615 65.710 26.935 ;
        RECT 66.040 26.615 66.300 26.935 ;
        RECT 66.830 26.615 67.090 26.935 ;
        RECT 65.465 25.365 65.695 26.615 ;
        RECT 66.055 25.365 66.285 26.615 ;
        RECT 66.845 25.365 67.075 26.615 ;
        RECT 67.315 25.160 67.575 25.665 ;
        RECT 64.225 24.930 65.415 25.160 ;
        RECT 66.335 24.930 67.575 25.160 ;
        RECT 68.000 24.715 68.355 26.905 ;
        RECT 63.400 24.440 64.065 24.715 ;
        RECT 67.685 24.440 68.355 24.715 ;
        RECT 63.400 22.335 63.755 24.440 ;
        RECT 64.175 24.015 65.415 24.245 ;
        RECT 66.335 24.015 67.525 24.245 ;
        RECT 64.175 23.590 64.435 24.015 ;
        RECT 64.675 22.575 64.905 23.810 ;
        RECT 65.465 22.575 65.695 23.810 ;
        RECT 66.055 22.575 66.285 23.810 ;
        RECT 56.655 21.205 56.915 21.995 ;
        RECT 53.515 20.975 54.755 21.205 ;
        RECT 55.675 20.975 56.915 21.205 ;
        RECT 58.840 21.205 59.100 22.085 ;
        RECT 59.340 21.365 59.570 22.255 ;
        RECT 60.130 21.365 60.360 22.255 ;
        RECT 60.720 21.365 60.950 22.255 ;
        RECT 61.510 21.365 61.740 22.330 ;
        RECT 64.660 22.255 64.920 22.575 ;
        RECT 65.450 22.255 65.710 22.575 ;
        RECT 66.040 22.255 66.300 22.575 ;
        RECT 66.845 22.500 67.075 23.810 ;
        RECT 67.265 22.940 67.525 24.015 ;
        RECT 67.685 22.500 67.855 24.440 ;
        RECT 66.845 22.330 67.855 22.500 ;
        RECT 68.000 22.330 68.355 24.440 ;
        RECT 68.725 24.715 69.080 26.910 ;
        RECT 70.000 26.845 70.230 27.810 ;
        RECT 70.790 26.935 71.020 27.810 ;
        RECT 71.380 26.935 71.610 27.810 ;
        RECT 72.170 26.935 72.400 27.810 ;
        RECT 72.640 27.180 72.900 27.970 ;
        RECT 74.835 27.970 76.075 28.200 ;
        RECT 76.995 27.970 78.235 28.200 ;
        RECT 74.835 27.275 75.095 27.970 ;
        RECT 69.220 26.675 70.230 26.845 ;
        RECT 69.220 24.715 69.390 26.675 ;
        RECT 69.550 25.160 69.810 26.295 ;
        RECT 70.000 25.365 70.230 26.675 ;
        RECT 70.775 26.615 71.035 26.935 ;
        RECT 71.365 26.615 71.625 26.935 ;
        RECT 72.155 26.615 72.415 26.935 ;
        RECT 70.790 25.365 71.020 26.615 ;
        RECT 71.380 25.365 71.610 26.615 ;
        RECT 72.170 25.365 72.400 26.615 ;
        RECT 72.640 25.160 72.900 25.665 ;
        RECT 69.550 24.930 70.740 25.160 ;
        RECT 71.660 24.930 72.900 25.160 ;
        RECT 73.325 24.715 73.680 26.905 ;
        RECT 68.725 24.440 69.390 24.715 ;
        RECT 73.010 24.440 73.680 24.715 ;
        RECT 68.725 22.335 69.080 24.440 ;
        RECT 69.500 24.015 70.740 24.245 ;
        RECT 71.660 24.015 72.850 24.245 ;
        RECT 69.500 23.590 69.760 24.015 ;
        RECT 70.000 22.575 70.230 23.810 ;
        RECT 70.790 22.575 71.020 23.810 ;
        RECT 71.380 22.575 71.610 23.810 ;
        RECT 61.980 21.205 62.240 21.995 ;
        RECT 58.840 20.975 60.080 21.205 ;
        RECT 61.000 20.975 62.240 21.205 ;
        RECT 64.175 21.205 64.435 22.085 ;
        RECT 64.675 21.365 64.905 22.255 ;
        RECT 65.465 21.365 65.695 22.255 ;
        RECT 66.055 21.365 66.285 22.255 ;
        RECT 66.845 21.365 67.075 22.330 ;
        RECT 69.985 22.255 70.245 22.575 ;
        RECT 70.775 22.255 71.035 22.575 ;
        RECT 71.365 22.255 71.625 22.575 ;
        RECT 72.170 22.500 72.400 23.810 ;
        RECT 72.590 22.940 72.850 24.015 ;
        RECT 73.010 22.500 73.180 24.440 ;
        RECT 72.170 22.330 73.180 22.500 ;
        RECT 73.325 22.330 73.680 24.440 ;
        RECT 74.060 24.715 74.415 26.910 ;
        RECT 75.335 26.845 75.565 27.810 ;
        RECT 76.125 26.935 76.355 27.810 ;
        RECT 76.715 26.935 76.945 27.810 ;
        RECT 77.505 26.935 77.735 27.810 ;
        RECT 77.975 27.180 78.235 27.970 ;
        RECT 80.160 27.970 81.400 28.200 ;
        RECT 82.320 27.970 83.560 28.200 ;
        RECT 80.160 27.275 80.420 27.970 ;
        RECT 74.555 26.675 75.565 26.845 ;
        RECT 74.555 24.715 74.725 26.675 ;
        RECT 74.885 25.160 75.145 26.295 ;
        RECT 75.335 25.365 75.565 26.675 ;
        RECT 76.110 26.615 76.370 26.935 ;
        RECT 76.700 26.615 76.960 26.935 ;
        RECT 77.490 26.615 77.750 26.935 ;
        RECT 76.125 25.365 76.355 26.615 ;
        RECT 76.715 25.365 76.945 26.615 ;
        RECT 77.505 25.365 77.735 26.615 ;
        RECT 77.975 25.160 78.235 25.665 ;
        RECT 74.885 24.930 76.075 25.160 ;
        RECT 76.995 24.930 78.235 25.160 ;
        RECT 78.660 24.715 79.015 26.905 ;
        RECT 74.060 24.440 74.725 24.715 ;
        RECT 78.345 24.440 79.015 24.715 ;
        RECT 74.060 22.335 74.415 24.440 ;
        RECT 74.835 24.015 76.075 24.245 ;
        RECT 76.995 24.015 78.185 24.245 ;
        RECT 74.835 23.590 75.095 24.015 ;
        RECT 75.335 22.575 75.565 23.810 ;
        RECT 76.125 22.575 76.355 23.810 ;
        RECT 76.715 22.575 76.945 23.810 ;
        RECT 67.315 21.205 67.575 21.995 ;
        RECT 64.175 20.975 65.415 21.205 ;
        RECT 66.335 20.975 67.575 21.205 ;
        RECT 69.500 21.205 69.760 22.085 ;
        RECT 70.000 21.365 70.230 22.255 ;
        RECT 70.790 21.365 71.020 22.255 ;
        RECT 71.380 21.365 71.610 22.255 ;
        RECT 72.170 21.365 72.400 22.330 ;
        RECT 75.320 22.255 75.580 22.575 ;
        RECT 76.110 22.255 76.370 22.575 ;
        RECT 76.700 22.255 76.960 22.575 ;
        RECT 77.505 22.500 77.735 23.810 ;
        RECT 77.925 22.940 78.185 24.015 ;
        RECT 78.345 22.500 78.515 24.440 ;
        RECT 77.505 22.330 78.515 22.500 ;
        RECT 78.660 22.330 79.015 24.440 ;
        RECT 79.385 24.715 79.740 26.910 ;
        RECT 80.660 26.845 80.890 27.810 ;
        RECT 81.450 26.935 81.680 27.810 ;
        RECT 82.040 26.935 82.270 27.810 ;
        RECT 82.830 26.935 83.060 27.810 ;
        RECT 83.300 27.180 83.560 27.970 ;
        RECT 85.495 27.970 86.735 28.200 ;
        RECT 87.655 27.970 88.895 28.200 ;
        RECT 85.495 27.275 85.755 27.970 ;
        RECT 79.880 26.675 80.890 26.845 ;
        RECT 79.880 24.715 80.050 26.675 ;
        RECT 80.210 25.160 80.470 26.295 ;
        RECT 80.660 25.365 80.890 26.675 ;
        RECT 81.435 26.615 81.695 26.935 ;
        RECT 82.025 26.615 82.285 26.935 ;
        RECT 82.815 26.615 83.075 26.935 ;
        RECT 81.450 25.365 81.680 26.615 ;
        RECT 82.040 25.365 82.270 26.615 ;
        RECT 82.830 25.365 83.060 26.615 ;
        RECT 83.300 25.160 83.560 25.665 ;
        RECT 80.210 24.930 81.400 25.160 ;
        RECT 82.320 24.930 83.560 25.160 ;
        RECT 83.985 24.715 84.340 26.905 ;
        RECT 79.385 24.440 80.050 24.715 ;
        RECT 83.670 24.440 84.340 24.715 ;
        RECT 79.385 22.335 79.740 24.440 ;
        RECT 80.160 24.015 81.400 24.245 ;
        RECT 82.320 24.015 83.510 24.245 ;
        RECT 80.160 23.590 80.420 24.015 ;
        RECT 80.660 22.575 80.890 23.810 ;
        RECT 81.450 22.575 81.680 23.810 ;
        RECT 82.040 22.575 82.270 23.810 ;
        RECT 72.640 21.205 72.900 21.995 ;
        RECT 69.500 20.975 70.740 21.205 ;
        RECT 71.660 20.975 72.900 21.205 ;
        RECT 74.835 21.205 75.095 22.085 ;
        RECT 75.335 21.365 75.565 22.255 ;
        RECT 76.125 21.365 76.355 22.255 ;
        RECT 76.715 21.365 76.945 22.255 ;
        RECT 77.505 21.365 77.735 22.330 ;
        RECT 80.645 22.255 80.905 22.575 ;
        RECT 81.435 22.255 81.695 22.575 ;
        RECT 82.025 22.255 82.285 22.575 ;
        RECT 82.830 22.500 83.060 23.810 ;
        RECT 83.250 22.940 83.510 24.015 ;
        RECT 83.670 22.500 83.840 24.440 ;
        RECT 82.830 22.330 83.840 22.500 ;
        RECT 83.985 22.330 84.340 24.440 ;
        RECT 84.720 24.715 85.075 26.910 ;
        RECT 85.995 26.845 86.225 27.810 ;
        RECT 86.785 26.935 87.015 27.810 ;
        RECT 87.375 26.935 87.605 27.810 ;
        RECT 88.165 26.935 88.395 27.810 ;
        RECT 88.635 27.180 88.895 27.970 ;
        RECT 90.820 27.970 92.060 28.200 ;
        RECT 92.980 27.970 94.220 28.200 ;
        RECT 90.820 27.275 91.080 27.970 ;
        RECT 85.215 26.675 86.225 26.845 ;
        RECT 85.215 24.715 85.385 26.675 ;
        RECT 85.545 25.160 85.805 26.295 ;
        RECT 85.995 25.365 86.225 26.675 ;
        RECT 86.770 26.615 87.030 26.935 ;
        RECT 87.360 26.615 87.620 26.935 ;
        RECT 88.150 26.615 88.410 26.935 ;
        RECT 86.785 25.365 87.015 26.615 ;
        RECT 87.375 25.365 87.605 26.615 ;
        RECT 88.165 25.365 88.395 26.615 ;
        RECT 88.635 25.160 88.895 25.665 ;
        RECT 85.545 24.930 86.735 25.160 ;
        RECT 87.655 24.930 88.895 25.160 ;
        RECT 89.320 24.715 89.675 26.905 ;
        RECT 84.720 24.440 85.385 24.715 ;
        RECT 89.005 24.440 89.675 24.715 ;
        RECT 84.720 22.335 85.075 24.440 ;
        RECT 85.495 24.015 86.735 24.245 ;
        RECT 87.655 24.015 88.845 24.245 ;
        RECT 85.495 23.590 85.755 24.015 ;
        RECT 85.995 22.575 86.225 23.810 ;
        RECT 86.785 22.575 87.015 23.810 ;
        RECT 87.375 22.575 87.605 23.810 ;
        RECT 77.975 21.205 78.235 21.995 ;
        RECT 74.835 20.975 76.075 21.205 ;
        RECT 76.995 20.975 78.235 21.205 ;
        RECT 80.160 21.205 80.420 22.085 ;
        RECT 80.660 21.365 80.890 22.255 ;
        RECT 81.450 21.365 81.680 22.255 ;
        RECT 82.040 21.365 82.270 22.255 ;
        RECT 82.830 21.365 83.060 22.330 ;
        RECT 85.980 22.255 86.240 22.575 ;
        RECT 86.770 22.255 87.030 22.575 ;
        RECT 87.360 22.255 87.620 22.575 ;
        RECT 88.165 22.500 88.395 23.810 ;
        RECT 88.585 22.940 88.845 24.015 ;
        RECT 89.005 22.500 89.175 24.440 ;
        RECT 88.165 22.330 89.175 22.500 ;
        RECT 89.320 22.330 89.675 24.440 ;
        RECT 90.045 24.715 90.400 26.910 ;
        RECT 91.320 26.845 91.550 27.810 ;
        RECT 92.110 26.935 92.340 27.810 ;
        RECT 92.700 26.935 92.930 27.810 ;
        RECT 93.490 26.935 93.720 27.810 ;
        RECT 93.960 27.180 94.220 27.970 ;
        RECT 96.155 27.970 97.395 28.200 ;
        RECT 98.315 27.970 99.555 28.200 ;
        RECT 96.155 27.275 96.415 27.970 ;
        RECT 90.540 26.675 91.550 26.845 ;
        RECT 90.540 24.715 90.710 26.675 ;
        RECT 90.870 25.160 91.130 26.295 ;
        RECT 91.320 25.365 91.550 26.675 ;
        RECT 92.095 26.615 92.355 26.935 ;
        RECT 92.685 26.615 92.945 26.935 ;
        RECT 93.475 26.615 93.735 26.935 ;
        RECT 92.110 25.365 92.340 26.615 ;
        RECT 92.700 25.365 92.930 26.615 ;
        RECT 93.490 25.365 93.720 26.615 ;
        RECT 93.960 25.160 94.220 25.665 ;
        RECT 90.870 24.930 92.060 25.160 ;
        RECT 92.980 24.930 94.220 25.160 ;
        RECT 94.645 24.715 95.000 26.905 ;
        RECT 90.045 24.440 90.710 24.715 ;
        RECT 94.330 24.440 95.000 24.715 ;
        RECT 90.045 22.335 90.400 24.440 ;
        RECT 90.820 24.015 92.060 24.245 ;
        RECT 92.980 24.015 94.170 24.245 ;
        RECT 90.820 23.590 91.080 24.015 ;
        RECT 91.320 22.575 91.550 23.810 ;
        RECT 92.110 22.575 92.340 23.810 ;
        RECT 92.700 22.575 92.930 23.810 ;
        RECT 83.300 21.205 83.560 21.995 ;
        RECT 80.160 20.975 81.400 21.205 ;
        RECT 82.320 20.975 83.560 21.205 ;
        RECT 85.495 21.205 85.755 22.085 ;
        RECT 85.995 21.365 86.225 22.255 ;
        RECT 86.785 21.365 87.015 22.255 ;
        RECT 87.375 21.365 87.605 22.255 ;
        RECT 88.165 21.365 88.395 22.330 ;
        RECT 91.305 22.255 91.565 22.575 ;
        RECT 92.095 22.255 92.355 22.575 ;
        RECT 92.685 22.255 92.945 22.575 ;
        RECT 93.490 22.500 93.720 23.810 ;
        RECT 93.910 22.940 94.170 24.015 ;
        RECT 94.330 22.500 94.500 24.440 ;
        RECT 93.490 22.330 94.500 22.500 ;
        RECT 94.645 22.330 95.000 24.440 ;
        RECT 95.380 24.715 95.735 26.910 ;
        RECT 96.655 26.845 96.885 27.810 ;
        RECT 97.445 26.935 97.675 27.810 ;
        RECT 98.035 26.935 98.265 27.810 ;
        RECT 98.825 26.935 99.055 27.810 ;
        RECT 99.295 27.180 99.555 27.970 ;
        RECT 101.480 27.970 102.720 28.200 ;
        RECT 103.640 27.970 104.880 28.200 ;
        RECT 101.480 27.275 101.740 27.970 ;
        RECT 95.875 26.675 96.885 26.845 ;
        RECT 95.875 24.715 96.045 26.675 ;
        RECT 96.205 25.160 96.465 26.295 ;
        RECT 96.655 25.365 96.885 26.675 ;
        RECT 97.430 26.615 97.690 26.935 ;
        RECT 98.020 26.615 98.280 26.935 ;
        RECT 98.810 26.615 99.070 26.935 ;
        RECT 97.445 25.365 97.675 26.615 ;
        RECT 98.035 25.365 98.265 26.615 ;
        RECT 98.825 25.365 99.055 26.615 ;
        RECT 99.295 25.160 99.555 25.665 ;
        RECT 96.205 24.930 97.395 25.160 ;
        RECT 98.315 24.930 99.555 25.160 ;
        RECT 99.980 24.715 100.335 26.905 ;
        RECT 95.380 24.440 96.045 24.715 ;
        RECT 99.665 24.440 100.335 24.715 ;
        RECT 95.380 22.335 95.735 24.440 ;
        RECT 96.155 24.015 97.395 24.245 ;
        RECT 98.315 24.015 99.505 24.245 ;
        RECT 96.155 23.590 96.415 24.015 ;
        RECT 96.655 22.575 96.885 23.810 ;
        RECT 97.445 22.575 97.675 23.810 ;
        RECT 98.035 22.575 98.265 23.810 ;
        RECT 88.635 21.205 88.895 21.995 ;
        RECT 85.495 20.975 86.735 21.205 ;
        RECT 87.655 20.975 88.895 21.205 ;
        RECT 90.820 21.205 91.080 22.085 ;
        RECT 91.320 21.365 91.550 22.255 ;
        RECT 92.110 21.365 92.340 22.255 ;
        RECT 92.700 21.365 92.930 22.255 ;
        RECT 93.490 21.365 93.720 22.330 ;
        RECT 96.640 22.255 96.900 22.575 ;
        RECT 97.430 22.255 97.690 22.575 ;
        RECT 98.020 22.255 98.280 22.575 ;
        RECT 98.825 22.500 99.055 23.810 ;
        RECT 99.245 22.940 99.505 24.015 ;
        RECT 99.665 22.500 99.835 24.440 ;
        RECT 98.825 22.330 99.835 22.500 ;
        RECT 99.980 22.330 100.335 24.440 ;
        RECT 100.705 24.715 101.060 26.910 ;
        RECT 101.980 26.845 102.210 27.810 ;
        RECT 102.770 26.935 103.000 27.810 ;
        RECT 103.360 26.935 103.590 27.810 ;
        RECT 104.150 26.935 104.380 27.810 ;
        RECT 104.620 27.180 104.880 27.970 ;
        RECT 106.815 27.970 108.055 28.200 ;
        RECT 108.975 27.970 110.215 28.200 ;
        RECT 106.815 27.275 107.075 27.970 ;
        RECT 101.200 26.675 102.210 26.845 ;
        RECT 101.200 24.715 101.370 26.675 ;
        RECT 101.530 25.160 101.790 26.295 ;
        RECT 101.980 25.365 102.210 26.675 ;
        RECT 102.755 26.615 103.015 26.935 ;
        RECT 103.345 26.615 103.605 26.935 ;
        RECT 104.135 26.615 104.395 26.935 ;
        RECT 102.770 25.365 103.000 26.615 ;
        RECT 103.360 25.365 103.590 26.615 ;
        RECT 104.150 25.365 104.380 26.615 ;
        RECT 104.620 25.160 104.880 25.665 ;
        RECT 101.530 24.930 102.720 25.160 ;
        RECT 103.640 24.930 104.880 25.160 ;
        RECT 105.305 24.715 105.660 26.905 ;
        RECT 100.705 24.440 101.370 24.715 ;
        RECT 104.990 24.440 105.660 24.715 ;
        RECT 100.705 22.335 101.060 24.440 ;
        RECT 101.480 24.015 102.720 24.245 ;
        RECT 103.640 24.015 104.830 24.245 ;
        RECT 101.480 23.590 101.740 24.015 ;
        RECT 101.980 22.575 102.210 23.810 ;
        RECT 102.770 22.575 103.000 23.810 ;
        RECT 103.360 22.575 103.590 23.810 ;
        RECT 93.960 21.205 94.220 21.995 ;
        RECT 90.820 20.975 92.060 21.205 ;
        RECT 92.980 20.975 94.220 21.205 ;
        RECT 96.155 21.205 96.415 22.085 ;
        RECT 96.655 21.365 96.885 22.255 ;
        RECT 97.445 21.365 97.675 22.255 ;
        RECT 98.035 21.365 98.265 22.255 ;
        RECT 98.825 21.365 99.055 22.330 ;
        RECT 101.965 22.255 102.225 22.575 ;
        RECT 102.755 22.255 103.015 22.575 ;
        RECT 103.345 22.255 103.605 22.575 ;
        RECT 104.150 22.500 104.380 23.810 ;
        RECT 104.570 22.940 104.830 24.015 ;
        RECT 104.990 22.500 105.160 24.440 ;
        RECT 104.150 22.330 105.160 22.500 ;
        RECT 105.305 22.330 105.660 24.440 ;
        RECT 106.040 24.715 106.395 26.910 ;
        RECT 107.315 26.845 107.545 27.810 ;
        RECT 108.105 26.935 108.335 27.810 ;
        RECT 108.695 26.935 108.925 27.810 ;
        RECT 109.485 26.935 109.715 27.810 ;
        RECT 109.955 27.180 110.215 27.970 ;
        RECT 112.140 27.970 113.380 28.200 ;
        RECT 114.300 27.970 115.540 28.200 ;
        RECT 112.140 27.275 112.400 27.970 ;
        RECT 106.535 26.675 107.545 26.845 ;
        RECT 106.535 24.715 106.705 26.675 ;
        RECT 106.865 25.160 107.125 26.295 ;
        RECT 107.315 25.365 107.545 26.675 ;
        RECT 108.090 26.615 108.350 26.935 ;
        RECT 108.680 26.615 108.940 26.935 ;
        RECT 109.470 26.615 109.730 26.935 ;
        RECT 108.105 25.365 108.335 26.615 ;
        RECT 108.695 25.365 108.925 26.615 ;
        RECT 109.485 25.365 109.715 26.615 ;
        RECT 109.955 25.160 110.215 25.665 ;
        RECT 106.865 24.930 108.055 25.160 ;
        RECT 108.975 24.930 110.215 25.160 ;
        RECT 110.640 24.715 110.995 26.905 ;
        RECT 106.040 24.440 106.705 24.715 ;
        RECT 110.325 24.440 110.995 24.715 ;
        RECT 106.040 22.335 106.395 24.440 ;
        RECT 106.815 24.015 108.055 24.245 ;
        RECT 108.975 24.015 110.165 24.245 ;
        RECT 106.815 23.590 107.075 24.015 ;
        RECT 107.315 22.575 107.545 23.810 ;
        RECT 108.105 22.575 108.335 23.810 ;
        RECT 108.695 22.575 108.925 23.810 ;
        RECT 99.295 21.205 99.555 21.995 ;
        RECT 96.155 20.975 97.395 21.205 ;
        RECT 98.315 20.975 99.555 21.205 ;
        RECT 101.480 21.205 101.740 22.085 ;
        RECT 101.980 21.365 102.210 22.255 ;
        RECT 102.770 21.365 103.000 22.255 ;
        RECT 103.360 21.365 103.590 22.255 ;
        RECT 104.150 21.365 104.380 22.330 ;
        RECT 107.300 22.255 107.560 22.575 ;
        RECT 108.090 22.255 108.350 22.575 ;
        RECT 108.680 22.255 108.940 22.575 ;
        RECT 109.485 22.500 109.715 23.810 ;
        RECT 109.905 22.940 110.165 24.015 ;
        RECT 110.325 22.500 110.495 24.440 ;
        RECT 109.485 22.330 110.495 22.500 ;
        RECT 110.640 22.330 110.995 24.440 ;
        RECT 111.365 24.715 111.720 26.910 ;
        RECT 112.640 26.845 112.870 27.810 ;
        RECT 113.430 26.935 113.660 27.810 ;
        RECT 114.020 26.935 114.250 27.810 ;
        RECT 114.810 26.935 115.040 27.810 ;
        RECT 115.280 27.180 115.540 27.970 ;
        RECT 117.475 27.970 118.715 28.200 ;
        RECT 119.635 27.970 120.875 28.200 ;
        RECT 117.475 27.275 117.735 27.970 ;
        RECT 111.860 26.675 112.870 26.845 ;
        RECT 111.860 24.715 112.030 26.675 ;
        RECT 112.190 25.160 112.450 26.295 ;
        RECT 112.640 25.365 112.870 26.675 ;
        RECT 113.415 26.615 113.675 26.935 ;
        RECT 114.005 26.615 114.265 26.935 ;
        RECT 114.795 26.615 115.055 26.935 ;
        RECT 113.430 25.365 113.660 26.615 ;
        RECT 114.020 25.365 114.250 26.615 ;
        RECT 114.810 25.365 115.040 26.615 ;
        RECT 115.280 25.160 115.540 25.665 ;
        RECT 112.190 24.930 113.380 25.160 ;
        RECT 114.300 24.930 115.540 25.160 ;
        RECT 115.965 24.715 116.320 26.905 ;
        RECT 111.365 24.440 112.030 24.715 ;
        RECT 115.650 24.440 116.320 24.715 ;
        RECT 111.365 22.335 111.720 24.440 ;
        RECT 112.140 24.015 113.380 24.245 ;
        RECT 114.300 24.015 115.490 24.245 ;
        RECT 112.140 23.590 112.400 24.015 ;
        RECT 112.640 22.575 112.870 23.810 ;
        RECT 113.430 22.575 113.660 23.810 ;
        RECT 114.020 22.575 114.250 23.810 ;
        RECT 104.620 21.205 104.880 21.995 ;
        RECT 101.480 20.975 102.720 21.205 ;
        RECT 103.640 20.975 104.880 21.205 ;
        RECT 106.815 21.205 107.075 22.085 ;
        RECT 107.315 21.365 107.545 22.255 ;
        RECT 108.105 21.365 108.335 22.255 ;
        RECT 108.695 21.365 108.925 22.255 ;
        RECT 109.485 21.365 109.715 22.330 ;
        RECT 112.625 22.255 112.885 22.575 ;
        RECT 113.415 22.255 113.675 22.575 ;
        RECT 114.005 22.255 114.265 22.575 ;
        RECT 114.810 22.500 115.040 23.810 ;
        RECT 115.230 22.940 115.490 24.015 ;
        RECT 115.650 22.500 115.820 24.440 ;
        RECT 114.810 22.330 115.820 22.500 ;
        RECT 115.965 22.330 116.320 24.440 ;
        RECT 116.700 24.715 117.055 26.910 ;
        RECT 117.975 26.845 118.205 27.810 ;
        RECT 118.765 26.935 118.995 27.810 ;
        RECT 119.355 26.935 119.585 27.810 ;
        RECT 120.145 26.935 120.375 27.810 ;
        RECT 120.615 27.180 120.875 27.970 ;
        RECT 117.195 26.675 118.205 26.845 ;
        RECT 117.195 24.715 117.365 26.675 ;
        RECT 117.525 25.160 117.785 26.295 ;
        RECT 117.975 25.365 118.205 26.675 ;
        RECT 118.750 26.615 119.010 26.935 ;
        RECT 119.340 26.615 119.600 26.935 ;
        RECT 120.130 26.615 120.390 26.935 ;
        RECT 118.765 25.365 118.995 26.615 ;
        RECT 119.355 25.365 119.585 26.615 ;
        RECT 120.145 25.365 120.375 26.615 ;
        RECT 120.615 25.160 120.875 25.665 ;
        RECT 117.525 24.930 118.715 25.160 ;
        RECT 119.635 24.930 120.875 25.160 ;
        RECT 121.300 24.715 121.655 26.905 ;
        RECT 116.700 24.440 117.365 24.715 ;
        RECT 120.985 24.440 121.655 24.715 ;
        RECT 116.700 22.335 117.055 24.440 ;
        RECT 117.475 24.015 118.715 24.245 ;
        RECT 119.635 24.015 120.825 24.245 ;
        RECT 117.475 23.590 117.735 24.015 ;
        RECT 117.975 22.575 118.205 23.810 ;
        RECT 118.765 22.575 118.995 23.810 ;
        RECT 119.355 22.575 119.585 23.810 ;
        RECT 109.955 21.205 110.215 21.995 ;
        RECT 106.815 20.975 108.055 21.205 ;
        RECT 108.975 20.975 110.215 21.205 ;
        RECT 112.140 21.205 112.400 22.085 ;
        RECT 112.640 21.365 112.870 22.255 ;
        RECT 113.430 21.365 113.660 22.255 ;
        RECT 114.020 21.365 114.250 22.255 ;
        RECT 114.810 21.365 115.040 22.330 ;
        RECT 117.960 22.255 118.220 22.575 ;
        RECT 118.750 22.255 119.010 22.575 ;
        RECT 119.340 22.255 119.600 22.575 ;
        RECT 120.145 22.500 120.375 23.810 ;
        RECT 120.565 22.940 120.825 24.015 ;
        RECT 120.985 22.500 121.155 24.440 ;
        RECT 120.145 22.330 121.155 22.500 ;
        RECT 121.300 22.330 121.655 24.440 ;
        RECT 122.025 24.715 122.380 26.925 ;
        RECT 123.300 26.845 123.530 27.810 ;
        RECT 124.090 26.935 124.320 27.810 ;
        RECT 124.680 26.935 124.910 27.810 ;
        RECT 125.470 26.935 125.700 27.810 ;
        RECT 122.520 26.675 123.530 26.845 ;
        RECT 122.520 24.715 122.690 26.675 ;
        RECT 123.300 25.365 123.530 26.675 ;
        RECT 124.075 26.615 124.335 26.935 ;
        RECT 124.665 26.615 124.925 26.935 ;
        RECT 125.455 26.615 125.715 26.935 ;
        RECT 124.090 25.365 124.320 26.615 ;
        RECT 124.680 25.365 124.910 26.615 ;
        RECT 125.470 25.365 125.700 26.615 ;
        RECT 126.625 24.715 126.980 26.925 ;
        RECT 122.025 24.440 122.690 24.715 ;
        RECT 126.310 24.440 126.980 24.715 ;
        RECT 122.025 22.350 122.380 24.440 ;
        RECT 123.300 22.575 123.530 23.810 ;
        RECT 124.090 22.575 124.320 23.810 ;
        RECT 124.680 22.575 124.910 23.810 ;
        RECT 115.280 21.205 115.540 21.995 ;
        RECT 112.140 20.975 113.380 21.205 ;
        RECT 114.300 20.975 115.540 21.205 ;
        RECT 117.475 21.205 117.735 22.085 ;
        RECT 117.975 21.365 118.205 22.255 ;
        RECT 118.765 21.365 118.995 22.255 ;
        RECT 119.355 21.365 119.585 22.255 ;
        RECT 120.145 21.365 120.375 22.330 ;
        RECT 123.285 22.255 123.545 22.575 ;
        RECT 124.075 22.255 124.335 22.575 ;
        RECT 124.665 22.255 124.925 22.575 ;
        RECT 125.470 22.500 125.700 23.810 ;
        RECT 126.310 22.500 126.480 24.440 ;
        RECT 125.470 22.330 126.480 22.500 ;
        RECT 126.625 22.350 126.980 24.440 ;
        RECT 120.615 21.205 120.875 21.995 ;
        RECT 123.300 21.365 123.530 22.255 ;
        RECT 124.090 21.365 124.320 22.255 ;
        RECT 124.680 21.365 124.910 22.255 ;
        RECT 125.470 21.365 125.700 22.330 ;
        RECT 117.475 20.975 118.715 21.205 ;
        RECT 119.635 20.975 120.875 21.205 ;
        RECT 37.520 20.435 38.760 20.665 ;
        RECT 39.680 20.435 40.920 20.665 ;
        RECT 10.500 19.910 10.820 20.395 ;
        RECT 16.115 20.020 26.850 20.255 ;
        RECT 10.500 19.580 11.960 19.910 ;
        RECT 10.500 19.360 10.820 19.580 ;
        RECT 12.400 18.835 12.720 19.825 ;
        RECT 14.585 19.580 16.005 19.905 ;
        RECT 19.990 19.450 26.850 20.020 ;
        RECT 16.115 19.215 26.850 19.450 ;
        RECT 12.425 18.820 12.715 18.835 ;
        RECT 27.665 17.435 27.925 17.440 ;
        RECT 25.540 16.835 27.985 17.435 ;
        RECT 10.510 15.315 10.810 16.765 ;
        RECT 15.985 16.600 27.985 16.835 ;
        RECT 11.745 16.215 13.345 16.505 ;
        RECT 14.165 16.215 20.945 16.450 ;
        RECT 21.425 16.400 27.985 16.600 ;
        RECT 31.420 17.180 31.775 19.390 ;
        RECT 32.695 19.310 32.925 20.275 ;
        RECT 33.485 19.400 33.715 20.275 ;
        RECT 34.075 19.400 34.305 20.275 ;
        RECT 34.865 19.400 35.095 20.275 ;
        RECT 37.520 19.740 37.780 20.435 ;
        RECT 31.915 19.140 32.925 19.310 ;
        RECT 31.915 17.180 32.085 19.140 ;
        RECT 32.695 17.830 32.925 19.140 ;
        RECT 33.470 19.080 33.730 19.400 ;
        RECT 34.060 19.080 34.320 19.400 ;
        RECT 34.850 19.080 35.110 19.400 ;
        RECT 33.485 17.830 33.715 19.080 ;
        RECT 34.075 17.830 34.305 19.080 ;
        RECT 34.865 17.830 35.095 19.080 ;
        RECT 36.020 17.180 36.375 19.390 ;
        RECT 31.420 16.905 32.085 17.180 ;
        RECT 35.705 16.905 36.375 17.180 ;
        RECT 16.040 16.030 17.645 16.060 ;
        RECT 21.425 16.030 26.675 16.400 ;
        RECT 15.985 15.800 26.675 16.030 ;
        RECT 15.985 15.795 22.260 15.800 ;
        RECT 16.040 15.770 17.645 15.795 ;
        RECT 31.420 14.815 31.775 16.905 ;
        RECT 32.695 15.040 32.925 16.275 ;
        RECT 33.485 15.040 33.715 16.275 ;
        RECT 34.075 15.040 34.305 16.275 ;
        RECT 32.680 14.720 32.940 15.040 ;
        RECT 33.470 14.720 33.730 15.040 ;
        RECT 34.060 14.720 34.320 15.040 ;
        RECT 34.865 14.965 35.095 16.275 ;
        RECT 35.705 14.965 35.875 16.905 ;
        RECT 34.865 14.795 35.875 14.965 ;
        RECT 36.020 14.815 36.375 16.905 ;
        RECT 36.745 17.180 37.100 19.375 ;
        RECT 38.020 19.310 38.250 20.275 ;
        RECT 38.810 19.400 39.040 20.275 ;
        RECT 39.400 19.400 39.630 20.275 ;
        RECT 40.190 19.400 40.420 20.275 ;
        RECT 40.660 19.645 40.920 20.435 ;
        RECT 42.855 20.435 44.095 20.665 ;
        RECT 45.015 20.435 46.255 20.665 ;
        RECT 42.855 19.740 43.115 20.435 ;
        RECT 37.240 19.140 38.250 19.310 ;
        RECT 37.240 17.180 37.410 19.140 ;
        RECT 37.570 17.625 37.830 18.760 ;
        RECT 38.020 17.830 38.250 19.140 ;
        RECT 38.795 19.080 39.055 19.400 ;
        RECT 39.385 19.080 39.645 19.400 ;
        RECT 40.175 19.080 40.435 19.400 ;
        RECT 38.810 17.830 39.040 19.080 ;
        RECT 39.400 17.830 39.630 19.080 ;
        RECT 40.190 17.830 40.420 19.080 ;
        RECT 40.660 17.625 40.920 18.130 ;
        RECT 37.570 17.395 38.760 17.625 ;
        RECT 39.680 17.395 40.920 17.625 ;
        RECT 41.345 17.180 41.700 19.370 ;
        RECT 36.745 16.905 37.410 17.180 ;
        RECT 41.030 16.905 41.700 17.180 ;
        RECT 36.745 14.800 37.100 16.905 ;
        RECT 37.520 16.480 38.760 16.710 ;
        RECT 39.680 16.480 40.870 16.710 ;
        RECT 37.520 16.055 37.780 16.480 ;
        RECT 38.020 15.040 38.250 16.275 ;
        RECT 38.810 15.040 39.040 16.275 ;
        RECT 39.400 15.040 39.630 16.275 ;
        RECT 32.695 13.830 32.925 14.720 ;
        RECT 33.485 13.830 33.715 14.720 ;
        RECT 34.075 13.830 34.305 14.720 ;
        RECT 34.865 13.830 35.095 14.795 ;
        RECT 38.005 14.720 38.265 15.040 ;
        RECT 38.795 14.720 39.055 15.040 ;
        RECT 39.385 14.720 39.645 15.040 ;
        RECT 40.190 14.965 40.420 16.275 ;
        RECT 40.610 15.405 40.870 16.480 ;
        RECT 41.030 14.965 41.200 16.905 ;
        RECT 40.190 14.795 41.200 14.965 ;
        RECT 41.345 14.795 41.700 16.905 ;
        RECT 42.080 17.180 42.435 19.375 ;
        RECT 43.355 19.310 43.585 20.275 ;
        RECT 44.145 19.400 44.375 20.275 ;
        RECT 44.735 19.400 44.965 20.275 ;
        RECT 45.525 19.400 45.755 20.275 ;
        RECT 45.995 19.645 46.255 20.435 ;
        RECT 48.180 20.435 49.420 20.665 ;
        RECT 50.340 20.435 51.580 20.665 ;
        RECT 48.180 19.740 48.440 20.435 ;
        RECT 42.575 19.140 43.585 19.310 ;
        RECT 42.575 17.180 42.745 19.140 ;
        RECT 42.905 17.625 43.165 18.760 ;
        RECT 43.355 17.830 43.585 19.140 ;
        RECT 44.130 19.080 44.390 19.400 ;
        RECT 44.720 19.080 44.980 19.400 ;
        RECT 45.510 19.080 45.770 19.400 ;
        RECT 44.145 17.830 44.375 19.080 ;
        RECT 44.735 17.830 44.965 19.080 ;
        RECT 45.525 17.830 45.755 19.080 ;
        RECT 45.995 17.625 46.255 18.130 ;
        RECT 42.905 17.395 44.095 17.625 ;
        RECT 45.015 17.395 46.255 17.625 ;
        RECT 46.680 17.180 47.035 19.370 ;
        RECT 42.080 16.905 42.745 17.180 ;
        RECT 46.365 16.905 47.035 17.180 ;
        RECT 42.080 14.800 42.435 16.905 ;
        RECT 42.855 16.480 44.095 16.710 ;
        RECT 45.015 16.480 46.205 16.710 ;
        RECT 42.855 16.055 43.115 16.480 ;
        RECT 43.355 15.040 43.585 16.275 ;
        RECT 44.145 15.040 44.375 16.275 ;
        RECT 44.735 15.040 44.965 16.275 ;
        RECT 37.520 13.670 37.780 14.550 ;
        RECT 38.020 13.830 38.250 14.720 ;
        RECT 38.810 13.830 39.040 14.720 ;
        RECT 39.400 13.830 39.630 14.720 ;
        RECT 40.190 13.830 40.420 14.795 ;
        RECT 43.340 14.720 43.600 15.040 ;
        RECT 44.130 14.720 44.390 15.040 ;
        RECT 44.720 14.720 44.980 15.040 ;
        RECT 45.525 14.965 45.755 16.275 ;
        RECT 45.945 15.405 46.205 16.480 ;
        RECT 46.365 14.965 46.535 16.905 ;
        RECT 45.525 14.795 46.535 14.965 ;
        RECT 46.680 14.795 47.035 16.905 ;
        RECT 47.405 17.180 47.760 19.375 ;
        RECT 48.680 19.310 48.910 20.275 ;
        RECT 49.470 19.400 49.700 20.275 ;
        RECT 50.060 19.400 50.290 20.275 ;
        RECT 50.850 19.400 51.080 20.275 ;
        RECT 51.320 19.645 51.580 20.435 ;
        RECT 53.515 20.435 54.755 20.665 ;
        RECT 55.675 20.435 56.915 20.665 ;
        RECT 53.515 19.740 53.775 20.435 ;
        RECT 47.900 19.140 48.910 19.310 ;
        RECT 47.900 17.180 48.070 19.140 ;
        RECT 48.230 17.625 48.490 18.760 ;
        RECT 48.680 17.830 48.910 19.140 ;
        RECT 49.455 19.080 49.715 19.400 ;
        RECT 50.045 19.080 50.305 19.400 ;
        RECT 50.835 19.080 51.095 19.400 ;
        RECT 49.470 17.830 49.700 19.080 ;
        RECT 50.060 17.830 50.290 19.080 ;
        RECT 50.850 17.830 51.080 19.080 ;
        RECT 51.320 17.625 51.580 18.130 ;
        RECT 48.230 17.395 49.420 17.625 ;
        RECT 50.340 17.395 51.580 17.625 ;
        RECT 52.005 17.180 52.360 19.370 ;
        RECT 47.405 16.905 48.070 17.180 ;
        RECT 51.690 16.905 52.360 17.180 ;
        RECT 47.405 14.800 47.760 16.905 ;
        RECT 48.180 16.480 49.420 16.710 ;
        RECT 50.340 16.480 51.530 16.710 ;
        RECT 48.180 16.055 48.440 16.480 ;
        RECT 48.680 15.040 48.910 16.275 ;
        RECT 49.470 15.040 49.700 16.275 ;
        RECT 50.060 15.040 50.290 16.275 ;
        RECT 40.660 13.670 40.920 14.460 ;
        RECT 37.520 13.440 38.760 13.670 ;
        RECT 39.680 13.440 40.920 13.670 ;
        RECT 42.855 13.670 43.115 14.550 ;
        RECT 43.355 13.830 43.585 14.720 ;
        RECT 44.145 13.830 44.375 14.720 ;
        RECT 44.735 13.830 44.965 14.720 ;
        RECT 45.525 13.830 45.755 14.795 ;
        RECT 48.665 14.720 48.925 15.040 ;
        RECT 49.455 14.720 49.715 15.040 ;
        RECT 50.045 14.720 50.305 15.040 ;
        RECT 50.850 14.965 51.080 16.275 ;
        RECT 51.270 15.405 51.530 16.480 ;
        RECT 51.690 14.965 51.860 16.905 ;
        RECT 50.850 14.795 51.860 14.965 ;
        RECT 52.005 14.795 52.360 16.905 ;
        RECT 52.740 17.180 53.095 19.375 ;
        RECT 54.015 19.310 54.245 20.275 ;
        RECT 54.805 19.400 55.035 20.275 ;
        RECT 55.395 19.400 55.625 20.275 ;
        RECT 56.185 19.400 56.415 20.275 ;
        RECT 56.655 19.645 56.915 20.435 ;
        RECT 58.840 20.435 60.080 20.665 ;
        RECT 61.000 20.435 62.240 20.665 ;
        RECT 58.840 19.740 59.100 20.435 ;
        RECT 53.235 19.140 54.245 19.310 ;
        RECT 53.235 17.180 53.405 19.140 ;
        RECT 53.565 17.625 53.825 18.760 ;
        RECT 54.015 17.830 54.245 19.140 ;
        RECT 54.790 19.080 55.050 19.400 ;
        RECT 55.380 19.080 55.640 19.400 ;
        RECT 56.170 19.080 56.430 19.400 ;
        RECT 54.805 17.830 55.035 19.080 ;
        RECT 55.395 17.830 55.625 19.080 ;
        RECT 56.185 17.830 56.415 19.080 ;
        RECT 56.655 17.625 56.915 18.130 ;
        RECT 53.565 17.395 54.755 17.625 ;
        RECT 55.675 17.395 56.915 17.625 ;
        RECT 57.340 17.180 57.695 19.370 ;
        RECT 52.740 16.905 53.405 17.180 ;
        RECT 57.025 16.905 57.695 17.180 ;
        RECT 52.740 14.800 53.095 16.905 ;
        RECT 53.515 16.480 54.755 16.710 ;
        RECT 55.675 16.480 56.865 16.710 ;
        RECT 53.515 16.055 53.775 16.480 ;
        RECT 54.015 15.040 54.245 16.275 ;
        RECT 54.805 15.040 55.035 16.275 ;
        RECT 55.395 15.040 55.625 16.275 ;
        RECT 45.995 13.670 46.255 14.460 ;
        RECT 42.855 13.440 44.095 13.670 ;
        RECT 45.015 13.440 46.255 13.670 ;
        RECT 48.180 13.670 48.440 14.550 ;
        RECT 48.680 13.830 48.910 14.720 ;
        RECT 49.470 13.830 49.700 14.720 ;
        RECT 50.060 13.830 50.290 14.720 ;
        RECT 50.850 13.830 51.080 14.795 ;
        RECT 54.000 14.720 54.260 15.040 ;
        RECT 54.790 14.720 55.050 15.040 ;
        RECT 55.380 14.720 55.640 15.040 ;
        RECT 56.185 14.965 56.415 16.275 ;
        RECT 56.605 15.405 56.865 16.480 ;
        RECT 57.025 14.965 57.195 16.905 ;
        RECT 56.185 14.795 57.195 14.965 ;
        RECT 57.340 14.795 57.695 16.905 ;
        RECT 58.065 17.180 58.420 19.375 ;
        RECT 59.340 19.310 59.570 20.275 ;
        RECT 60.130 19.400 60.360 20.275 ;
        RECT 60.720 19.400 60.950 20.275 ;
        RECT 61.510 19.400 61.740 20.275 ;
        RECT 61.980 19.645 62.240 20.435 ;
        RECT 64.175 20.435 65.415 20.665 ;
        RECT 66.335 20.435 67.575 20.665 ;
        RECT 64.175 19.740 64.435 20.435 ;
        RECT 58.560 19.140 59.570 19.310 ;
        RECT 58.560 17.180 58.730 19.140 ;
        RECT 58.890 17.625 59.150 18.760 ;
        RECT 59.340 17.830 59.570 19.140 ;
        RECT 60.115 19.080 60.375 19.400 ;
        RECT 60.705 19.080 60.965 19.400 ;
        RECT 61.495 19.080 61.755 19.400 ;
        RECT 60.130 17.830 60.360 19.080 ;
        RECT 60.720 17.830 60.950 19.080 ;
        RECT 61.510 17.830 61.740 19.080 ;
        RECT 61.980 17.625 62.240 18.130 ;
        RECT 58.890 17.395 60.080 17.625 ;
        RECT 61.000 17.395 62.240 17.625 ;
        RECT 62.665 17.180 63.020 19.370 ;
        RECT 58.065 16.905 58.730 17.180 ;
        RECT 62.350 16.905 63.020 17.180 ;
        RECT 58.065 14.800 58.420 16.905 ;
        RECT 58.840 16.480 60.080 16.710 ;
        RECT 61.000 16.480 62.190 16.710 ;
        RECT 58.840 16.055 59.100 16.480 ;
        RECT 59.340 15.040 59.570 16.275 ;
        RECT 60.130 15.040 60.360 16.275 ;
        RECT 60.720 15.040 60.950 16.275 ;
        RECT 51.320 13.670 51.580 14.460 ;
        RECT 48.180 13.440 49.420 13.670 ;
        RECT 50.340 13.440 51.580 13.670 ;
        RECT 53.515 13.670 53.775 14.550 ;
        RECT 54.015 13.830 54.245 14.720 ;
        RECT 54.805 13.830 55.035 14.720 ;
        RECT 55.395 13.830 55.625 14.720 ;
        RECT 56.185 13.830 56.415 14.795 ;
        RECT 59.325 14.720 59.585 15.040 ;
        RECT 60.115 14.720 60.375 15.040 ;
        RECT 60.705 14.720 60.965 15.040 ;
        RECT 61.510 14.965 61.740 16.275 ;
        RECT 61.930 15.405 62.190 16.480 ;
        RECT 62.350 14.965 62.520 16.905 ;
        RECT 61.510 14.795 62.520 14.965 ;
        RECT 62.665 14.795 63.020 16.905 ;
        RECT 63.400 17.180 63.755 19.375 ;
        RECT 64.675 19.310 64.905 20.275 ;
        RECT 65.465 19.400 65.695 20.275 ;
        RECT 66.055 19.400 66.285 20.275 ;
        RECT 66.845 19.400 67.075 20.275 ;
        RECT 67.315 19.645 67.575 20.435 ;
        RECT 69.500 20.435 70.740 20.665 ;
        RECT 71.660 20.435 72.900 20.665 ;
        RECT 69.500 19.740 69.760 20.435 ;
        RECT 63.895 19.140 64.905 19.310 ;
        RECT 63.895 17.180 64.065 19.140 ;
        RECT 64.225 17.625 64.485 18.760 ;
        RECT 64.675 17.830 64.905 19.140 ;
        RECT 65.450 19.080 65.710 19.400 ;
        RECT 66.040 19.080 66.300 19.400 ;
        RECT 66.830 19.080 67.090 19.400 ;
        RECT 65.465 17.830 65.695 19.080 ;
        RECT 66.055 17.830 66.285 19.080 ;
        RECT 66.845 17.830 67.075 19.080 ;
        RECT 67.315 17.625 67.575 18.130 ;
        RECT 64.225 17.395 65.415 17.625 ;
        RECT 66.335 17.395 67.575 17.625 ;
        RECT 68.000 17.180 68.355 19.370 ;
        RECT 63.400 16.905 64.065 17.180 ;
        RECT 67.685 16.905 68.355 17.180 ;
        RECT 63.400 14.800 63.755 16.905 ;
        RECT 64.175 16.480 65.415 16.710 ;
        RECT 66.335 16.480 67.525 16.710 ;
        RECT 64.175 16.055 64.435 16.480 ;
        RECT 64.675 15.040 64.905 16.275 ;
        RECT 65.465 15.040 65.695 16.275 ;
        RECT 66.055 15.040 66.285 16.275 ;
        RECT 56.655 13.670 56.915 14.460 ;
        RECT 53.515 13.440 54.755 13.670 ;
        RECT 55.675 13.440 56.915 13.670 ;
        RECT 58.840 13.670 59.100 14.550 ;
        RECT 59.340 13.830 59.570 14.720 ;
        RECT 60.130 13.830 60.360 14.720 ;
        RECT 60.720 13.830 60.950 14.720 ;
        RECT 61.510 13.830 61.740 14.795 ;
        RECT 64.660 14.720 64.920 15.040 ;
        RECT 65.450 14.720 65.710 15.040 ;
        RECT 66.040 14.720 66.300 15.040 ;
        RECT 66.845 14.965 67.075 16.275 ;
        RECT 67.265 15.405 67.525 16.480 ;
        RECT 67.685 14.965 67.855 16.905 ;
        RECT 66.845 14.795 67.855 14.965 ;
        RECT 68.000 14.795 68.355 16.905 ;
        RECT 68.725 17.180 69.080 19.375 ;
        RECT 70.000 19.310 70.230 20.275 ;
        RECT 70.790 19.400 71.020 20.275 ;
        RECT 71.380 19.400 71.610 20.275 ;
        RECT 72.170 19.400 72.400 20.275 ;
        RECT 72.640 19.645 72.900 20.435 ;
        RECT 74.835 20.435 76.075 20.665 ;
        RECT 76.995 20.435 78.235 20.665 ;
        RECT 74.835 19.740 75.095 20.435 ;
        RECT 69.220 19.140 70.230 19.310 ;
        RECT 69.220 17.180 69.390 19.140 ;
        RECT 69.550 17.625 69.810 18.760 ;
        RECT 70.000 17.830 70.230 19.140 ;
        RECT 70.775 19.080 71.035 19.400 ;
        RECT 71.365 19.080 71.625 19.400 ;
        RECT 72.155 19.080 72.415 19.400 ;
        RECT 70.790 17.830 71.020 19.080 ;
        RECT 71.380 17.830 71.610 19.080 ;
        RECT 72.170 17.830 72.400 19.080 ;
        RECT 72.640 17.625 72.900 18.130 ;
        RECT 69.550 17.395 70.740 17.625 ;
        RECT 71.660 17.395 72.900 17.625 ;
        RECT 73.325 17.180 73.680 19.370 ;
        RECT 68.725 16.905 69.390 17.180 ;
        RECT 73.010 16.905 73.680 17.180 ;
        RECT 68.725 14.800 69.080 16.905 ;
        RECT 69.500 16.480 70.740 16.710 ;
        RECT 71.660 16.480 72.850 16.710 ;
        RECT 69.500 16.055 69.760 16.480 ;
        RECT 70.000 15.040 70.230 16.275 ;
        RECT 70.790 15.040 71.020 16.275 ;
        RECT 71.380 15.040 71.610 16.275 ;
        RECT 61.980 13.670 62.240 14.460 ;
        RECT 58.840 13.440 60.080 13.670 ;
        RECT 61.000 13.440 62.240 13.670 ;
        RECT 64.175 13.670 64.435 14.550 ;
        RECT 64.675 13.830 64.905 14.720 ;
        RECT 65.465 13.830 65.695 14.720 ;
        RECT 66.055 13.830 66.285 14.720 ;
        RECT 66.845 13.830 67.075 14.795 ;
        RECT 69.985 14.720 70.245 15.040 ;
        RECT 70.775 14.720 71.035 15.040 ;
        RECT 71.365 14.720 71.625 15.040 ;
        RECT 72.170 14.965 72.400 16.275 ;
        RECT 72.590 15.405 72.850 16.480 ;
        RECT 73.010 14.965 73.180 16.905 ;
        RECT 72.170 14.795 73.180 14.965 ;
        RECT 73.325 14.795 73.680 16.905 ;
        RECT 74.060 17.180 74.415 19.375 ;
        RECT 75.335 19.310 75.565 20.275 ;
        RECT 76.125 19.400 76.355 20.275 ;
        RECT 76.715 19.400 76.945 20.275 ;
        RECT 77.505 19.400 77.735 20.275 ;
        RECT 77.975 19.645 78.235 20.435 ;
        RECT 80.160 20.435 81.400 20.665 ;
        RECT 82.320 20.435 83.560 20.665 ;
        RECT 80.160 19.740 80.420 20.435 ;
        RECT 74.555 19.140 75.565 19.310 ;
        RECT 74.555 17.180 74.725 19.140 ;
        RECT 74.885 17.625 75.145 18.760 ;
        RECT 75.335 17.830 75.565 19.140 ;
        RECT 76.110 19.080 76.370 19.400 ;
        RECT 76.700 19.080 76.960 19.400 ;
        RECT 77.490 19.080 77.750 19.400 ;
        RECT 76.125 17.830 76.355 19.080 ;
        RECT 76.715 17.830 76.945 19.080 ;
        RECT 77.505 17.830 77.735 19.080 ;
        RECT 77.975 17.625 78.235 18.130 ;
        RECT 74.885 17.395 76.075 17.625 ;
        RECT 76.995 17.395 78.235 17.625 ;
        RECT 78.660 17.180 79.015 19.370 ;
        RECT 74.060 16.905 74.725 17.180 ;
        RECT 78.345 16.905 79.015 17.180 ;
        RECT 74.060 14.800 74.415 16.905 ;
        RECT 74.835 16.480 76.075 16.710 ;
        RECT 76.995 16.480 78.185 16.710 ;
        RECT 74.835 16.055 75.095 16.480 ;
        RECT 75.335 15.040 75.565 16.275 ;
        RECT 76.125 15.040 76.355 16.275 ;
        RECT 76.715 15.040 76.945 16.275 ;
        RECT 67.315 13.670 67.575 14.460 ;
        RECT 64.175 13.440 65.415 13.670 ;
        RECT 66.335 13.440 67.575 13.670 ;
        RECT 69.500 13.670 69.760 14.550 ;
        RECT 70.000 13.830 70.230 14.720 ;
        RECT 70.790 13.830 71.020 14.720 ;
        RECT 71.380 13.830 71.610 14.720 ;
        RECT 72.170 13.830 72.400 14.795 ;
        RECT 75.320 14.720 75.580 15.040 ;
        RECT 76.110 14.720 76.370 15.040 ;
        RECT 76.700 14.720 76.960 15.040 ;
        RECT 77.505 14.965 77.735 16.275 ;
        RECT 77.925 15.405 78.185 16.480 ;
        RECT 78.345 14.965 78.515 16.905 ;
        RECT 77.505 14.795 78.515 14.965 ;
        RECT 78.660 14.795 79.015 16.905 ;
        RECT 79.385 17.180 79.740 19.375 ;
        RECT 80.660 19.310 80.890 20.275 ;
        RECT 81.450 19.400 81.680 20.275 ;
        RECT 82.040 19.400 82.270 20.275 ;
        RECT 82.830 19.400 83.060 20.275 ;
        RECT 83.300 19.645 83.560 20.435 ;
        RECT 85.495 20.435 86.735 20.665 ;
        RECT 87.655 20.435 88.895 20.665 ;
        RECT 85.495 19.740 85.755 20.435 ;
        RECT 79.880 19.140 80.890 19.310 ;
        RECT 79.880 17.180 80.050 19.140 ;
        RECT 80.210 17.625 80.470 18.760 ;
        RECT 80.660 17.830 80.890 19.140 ;
        RECT 81.435 19.080 81.695 19.400 ;
        RECT 82.025 19.080 82.285 19.400 ;
        RECT 82.815 19.080 83.075 19.400 ;
        RECT 81.450 17.830 81.680 19.080 ;
        RECT 82.040 17.830 82.270 19.080 ;
        RECT 82.830 17.830 83.060 19.080 ;
        RECT 83.300 17.625 83.560 18.130 ;
        RECT 80.210 17.395 81.400 17.625 ;
        RECT 82.320 17.395 83.560 17.625 ;
        RECT 83.985 17.180 84.340 19.370 ;
        RECT 79.385 16.905 80.050 17.180 ;
        RECT 83.670 16.905 84.340 17.180 ;
        RECT 79.385 14.800 79.740 16.905 ;
        RECT 80.160 16.480 81.400 16.710 ;
        RECT 82.320 16.480 83.510 16.710 ;
        RECT 80.160 16.055 80.420 16.480 ;
        RECT 80.660 15.040 80.890 16.275 ;
        RECT 81.450 15.040 81.680 16.275 ;
        RECT 82.040 15.040 82.270 16.275 ;
        RECT 72.640 13.670 72.900 14.460 ;
        RECT 69.500 13.440 70.740 13.670 ;
        RECT 71.660 13.440 72.900 13.670 ;
        RECT 74.835 13.670 75.095 14.550 ;
        RECT 75.335 13.830 75.565 14.720 ;
        RECT 76.125 13.830 76.355 14.720 ;
        RECT 76.715 13.830 76.945 14.720 ;
        RECT 77.505 13.830 77.735 14.795 ;
        RECT 80.645 14.720 80.905 15.040 ;
        RECT 81.435 14.720 81.695 15.040 ;
        RECT 82.025 14.720 82.285 15.040 ;
        RECT 82.830 14.965 83.060 16.275 ;
        RECT 83.250 15.405 83.510 16.480 ;
        RECT 83.670 14.965 83.840 16.905 ;
        RECT 82.830 14.795 83.840 14.965 ;
        RECT 83.985 14.795 84.340 16.905 ;
        RECT 84.720 17.180 85.075 19.375 ;
        RECT 85.995 19.310 86.225 20.275 ;
        RECT 86.785 19.400 87.015 20.275 ;
        RECT 87.375 19.400 87.605 20.275 ;
        RECT 88.165 19.400 88.395 20.275 ;
        RECT 88.635 19.645 88.895 20.435 ;
        RECT 90.820 20.435 92.060 20.665 ;
        RECT 92.980 20.435 94.220 20.665 ;
        RECT 90.820 19.740 91.080 20.435 ;
        RECT 85.215 19.140 86.225 19.310 ;
        RECT 85.215 17.180 85.385 19.140 ;
        RECT 85.545 17.625 85.805 18.760 ;
        RECT 85.995 17.830 86.225 19.140 ;
        RECT 86.770 19.080 87.030 19.400 ;
        RECT 87.360 19.080 87.620 19.400 ;
        RECT 88.150 19.080 88.410 19.400 ;
        RECT 86.785 17.830 87.015 19.080 ;
        RECT 87.375 17.830 87.605 19.080 ;
        RECT 88.165 17.830 88.395 19.080 ;
        RECT 88.635 17.625 88.895 18.130 ;
        RECT 85.545 17.395 86.735 17.625 ;
        RECT 87.655 17.395 88.895 17.625 ;
        RECT 89.320 17.180 89.675 19.370 ;
        RECT 84.720 16.905 85.385 17.180 ;
        RECT 89.005 16.905 89.675 17.180 ;
        RECT 84.720 14.800 85.075 16.905 ;
        RECT 85.495 16.480 86.735 16.710 ;
        RECT 87.655 16.480 88.845 16.710 ;
        RECT 85.495 16.055 85.755 16.480 ;
        RECT 85.995 15.040 86.225 16.275 ;
        RECT 86.785 15.040 87.015 16.275 ;
        RECT 87.375 15.040 87.605 16.275 ;
        RECT 77.975 13.670 78.235 14.460 ;
        RECT 74.835 13.440 76.075 13.670 ;
        RECT 76.995 13.440 78.235 13.670 ;
        RECT 80.160 13.670 80.420 14.550 ;
        RECT 80.660 13.830 80.890 14.720 ;
        RECT 81.450 13.830 81.680 14.720 ;
        RECT 82.040 13.830 82.270 14.720 ;
        RECT 82.830 13.830 83.060 14.795 ;
        RECT 85.980 14.720 86.240 15.040 ;
        RECT 86.770 14.720 87.030 15.040 ;
        RECT 87.360 14.720 87.620 15.040 ;
        RECT 88.165 14.965 88.395 16.275 ;
        RECT 88.585 15.405 88.845 16.480 ;
        RECT 89.005 14.965 89.175 16.905 ;
        RECT 88.165 14.795 89.175 14.965 ;
        RECT 89.320 14.795 89.675 16.905 ;
        RECT 90.045 17.180 90.400 19.375 ;
        RECT 91.320 19.310 91.550 20.275 ;
        RECT 92.110 19.400 92.340 20.275 ;
        RECT 92.700 19.400 92.930 20.275 ;
        RECT 93.490 19.400 93.720 20.275 ;
        RECT 93.960 19.645 94.220 20.435 ;
        RECT 96.155 20.435 97.395 20.665 ;
        RECT 98.315 20.435 99.555 20.665 ;
        RECT 96.155 19.740 96.415 20.435 ;
        RECT 90.540 19.140 91.550 19.310 ;
        RECT 90.540 17.180 90.710 19.140 ;
        RECT 90.870 17.625 91.130 18.760 ;
        RECT 91.320 17.830 91.550 19.140 ;
        RECT 92.095 19.080 92.355 19.400 ;
        RECT 92.685 19.080 92.945 19.400 ;
        RECT 93.475 19.080 93.735 19.400 ;
        RECT 92.110 17.830 92.340 19.080 ;
        RECT 92.700 17.830 92.930 19.080 ;
        RECT 93.490 17.830 93.720 19.080 ;
        RECT 93.960 17.625 94.220 18.130 ;
        RECT 90.870 17.395 92.060 17.625 ;
        RECT 92.980 17.395 94.220 17.625 ;
        RECT 94.645 17.180 95.000 19.370 ;
        RECT 90.045 16.905 90.710 17.180 ;
        RECT 94.330 16.905 95.000 17.180 ;
        RECT 90.045 14.800 90.400 16.905 ;
        RECT 90.820 16.480 92.060 16.710 ;
        RECT 92.980 16.480 94.170 16.710 ;
        RECT 90.820 16.055 91.080 16.480 ;
        RECT 91.320 15.040 91.550 16.275 ;
        RECT 92.110 15.040 92.340 16.275 ;
        RECT 92.700 15.040 92.930 16.275 ;
        RECT 83.300 13.670 83.560 14.460 ;
        RECT 80.160 13.440 81.400 13.670 ;
        RECT 82.320 13.440 83.560 13.670 ;
        RECT 85.495 13.670 85.755 14.550 ;
        RECT 85.995 13.830 86.225 14.720 ;
        RECT 86.785 13.830 87.015 14.720 ;
        RECT 87.375 13.830 87.605 14.720 ;
        RECT 88.165 13.830 88.395 14.795 ;
        RECT 91.305 14.720 91.565 15.040 ;
        RECT 92.095 14.720 92.355 15.040 ;
        RECT 92.685 14.720 92.945 15.040 ;
        RECT 93.490 14.965 93.720 16.275 ;
        RECT 93.910 15.405 94.170 16.480 ;
        RECT 94.330 14.965 94.500 16.905 ;
        RECT 93.490 14.795 94.500 14.965 ;
        RECT 94.645 14.795 95.000 16.905 ;
        RECT 95.380 17.180 95.735 19.375 ;
        RECT 96.655 19.310 96.885 20.275 ;
        RECT 97.445 19.400 97.675 20.275 ;
        RECT 98.035 19.400 98.265 20.275 ;
        RECT 98.825 19.400 99.055 20.275 ;
        RECT 99.295 19.645 99.555 20.435 ;
        RECT 101.480 20.435 102.720 20.665 ;
        RECT 103.640 20.435 104.880 20.665 ;
        RECT 101.480 19.740 101.740 20.435 ;
        RECT 95.875 19.140 96.885 19.310 ;
        RECT 95.875 17.180 96.045 19.140 ;
        RECT 96.205 17.625 96.465 18.760 ;
        RECT 96.655 17.830 96.885 19.140 ;
        RECT 97.430 19.080 97.690 19.400 ;
        RECT 98.020 19.080 98.280 19.400 ;
        RECT 98.810 19.080 99.070 19.400 ;
        RECT 97.445 17.830 97.675 19.080 ;
        RECT 98.035 17.830 98.265 19.080 ;
        RECT 98.825 17.830 99.055 19.080 ;
        RECT 99.295 17.625 99.555 18.130 ;
        RECT 96.205 17.395 97.395 17.625 ;
        RECT 98.315 17.395 99.555 17.625 ;
        RECT 99.980 17.180 100.335 19.370 ;
        RECT 95.380 16.905 96.045 17.180 ;
        RECT 99.665 16.905 100.335 17.180 ;
        RECT 95.380 14.800 95.735 16.905 ;
        RECT 96.155 16.480 97.395 16.710 ;
        RECT 98.315 16.480 99.505 16.710 ;
        RECT 96.155 16.055 96.415 16.480 ;
        RECT 96.655 15.040 96.885 16.275 ;
        RECT 97.445 15.040 97.675 16.275 ;
        RECT 98.035 15.040 98.265 16.275 ;
        RECT 88.635 13.670 88.895 14.460 ;
        RECT 85.495 13.440 86.735 13.670 ;
        RECT 87.655 13.440 88.895 13.670 ;
        RECT 90.820 13.670 91.080 14.550 ;
        RECT 91.320 13.830 91.550 14.720 ;
        RECT 92.110 13.830 92.340 14.720 ;
        RECT 92.700 13.830 92.930 14.720 ;
        RECT 93.490 13.830 93.720 14.795 ;
        RECT 96.640 14.720 96.900 15.040 ;
        RECT 97.430 14.720 97.690 15.040 ;
        RECT 98.020 14.720 98.280 15.040 ;
        RECT 98.825 14.965 99.055 16.275 ;
        RECT 99.245 15.405 99.505 16.480 ;
        RECT 99.665 14.965 99.835 16.905 ;
        RECT 98.825 14.795 99.835 14.965 ;
        RECT 99.980 14.795 100.335 16.905 ;
        RECT 100.705 17.180 101.060 19.375 ;
        RECT 101.980 19.310 102.210 20.275 ;
        RECT 102.770 19.400 103.000 20.275 ;
        RECT 103.360 19.400 103.590 20.275 ;
        RECT 104.150 19.400 104.380 20.275 ;
        RECT 104.620 19.645 104.880 20.435 ;
        RECT 106.815 20.435 108.055 20.665 ;
        RECT 108.975 20.435 110.215 20.665 ;
        RECT 106.815 19.740 107.075 20.435 ;
        RECT 101.200 19.140 102.210 19.310 ;
        RECT 101.200 17.180 101.370 19.140 ;
        RECT 101.530 17.625 101.790 18.760 ;
        RECT 101.980 17.830 102.210 19.140 ;
        RECT 102.755 19.080 103.015 19.400 ;
        RECT 103.345 19.080 103.605 19.400 ;
        RECT 104.135 19.080 104.395 19.400 ;
        RECT 102.770 17.830 103.000 19.080 ;
        RECT 103.360 17.830 103.590 19.080 ;
        RECT 104.150 17.830 104.380 19.080 ;
        RECT 104.620 17.625 104.880 18.130 ;
        RECT 101.530 17.395 102.720 17.625 ;
        RECT 103.640 17.395 104.880 17.625 ;
        RECT 105.305 17.180 105.660 19.370 ;
        RECT 100.705 16.905 101.370 17.180 ;
        RECT 104.990 16.905 105.660 17.180 ;
        RECT 100.705 14.800 101.060 16.905 ;
        RECT 101.480 16.480 102.720 16.710 ;
        RECT 103.640 16.480 104.830 16.710 ;
        RECT 101.480 16.055 101.740 16.480 ;
        RECT 101.980 15.040 102.210 16.275 ;
        RECT 102.770 15.040 103.000 16.275 ;
        RECT 103.360 15.040 103.590 16.275 ;
        RECT 93.960 13.670 94.220 14.460 ;
        RECT 90.820 13.440 92.060 13.670 ;
        RECT 92.980 13.440 94.220 13.670 ;
        RECT 96.155 13.670 96.415 14.550 ;
        RECT 96.655 13.830 96.885 14.720 ;
        RECT 97.445 13.830 97.675 14.720 ;
        RECT 98.035 13.830 98.265 14.720 ;
        RECT 98.825 13.830 99.055 14.795 ;
        RECT 101.965 14.720 102.225 15.040 ;
        RECT 102.755 14.720 103.015 15.040 ;
        RECT 103.345 14.720 103.605 15.040 ;
        RECT 104.150 14.965 104.380 16.275 ;
        RECT 104.570 15.405 104.830 16.480 ;
        RECT 104.990 14.965 105.160 16.905 ;
        RECT 104.150 14.795 105.160 14.965 ;
        RECT 105.305 14.795 105.660 16.905 ;
        RECT 106.040 17.180 106.395 19.375 ;
        RECT 107.315 19.310 107.545 20.275 ;
        RECT 108.105 19.400 108.335 20.275 ;
        RECT 108.695 19.400 108.925 20.275 ;
        RECT 109.485 19.400 109.715 20.275 ;
        RECT 109.955 19.645 110.215 20.435 ;
        RECT 112.140 20.435 113.380 20.665 ;
        RECT 114.300 20.435 115.540 20.665 ;
        RECT 112.140 19.740 112.400 20.435 ;
        RECT 106.535 19.140 107.545 19.310 ;
        RECT 106.535 17.180 106.705 19.140 ;
        RECT 106.865 17.625 107.125 18.760 ;
        RECT 107.315 17.830 107.545 19.140 ;
        RECT 108.090 19.080 108.350 19.400 ;
        RECT 108.680 19.080 108.940 19.400 ;
        RECT 109.470 19.080 109.730 19.400 ;
        RECT 108.105 17.830 108.335 19.080 ;
        RECT 108.695 17.830 108.925 19.080 ;
        RECT 109.485 17.830 109.715 19.080 ;
        RECT 109.955 17.625 110.215 18.130 ;
        RECT 106.865 17.395 108.055 17.625 ;
        RECT 108.975 17.395 110.215 17.625 ;
        RECT 110.640 17.180 110.995 19.370 ;
        RECT 106.040 16.905 106.705 17.180 ;
        RECT 110.325 16.905 110.995 17.180 ;
        RECT 106.040 14.800 106.395 16.905 ;
        RECT 106.815 16.480 108.055 16.710 ;
        RECT 108.975 16.480 110.165 16.710 ;
        RECT 106.815 16.055 107.075 16.480 ;
        RECT 107.315 15.040 107.545 16.275 ;
        RECT 108.105 15.040 108.335 16.275 ;
        RECT 108.695 15.040 108.925 16.275 ;
        RECT 99.295 13.670 99.555 14.460 ;
        RECT 96.155 13.440 97.395 13.670 ;
        RECT 98.315 13.440 99.555 13.670 ;
        RECT 101.480 13.670 101.740 14.550 ;
        RECT 101.980 13.830 102.210 14.720 ;
        RECT 102.770 13.830 103.000 14.720 ;
        RECT 103.360 13.830 103.590 14.720 ;
        RECT 104.150 13.830 104.380 14.795 ;
        RECT 107.300 14.720 107.560 15.040 ;
        RECT 108.090 14.720 108.350 15.040 ;
        RECT 108.680 14.720 108.940 15.040 ;
        RECT 109.485 14.965 109.715 16.275 ;
        RECT 109.905 15.405 110.165 16.480 ;
        RECT 110.325 14.965 110.495 16.905 ;
        RECT 109.485 14.795 110.495 14.965 ;
        RECT 110.640 14.795 110.995 16.905 ;
        RECT 111.365 17.180 111.720 19.375 ;
        RECT 112.640 19.310 112.870 20.275 ;
        RECT 113.430 19.400 113.660 20.275 ;
        RECT 114.020 19.400 114.250 20.275 ;
        RECT 114.810 19.400 115.040 20.275 ;
        RECT 115.280 19.645 115.540 20.435 ;
        RECT 117.475 20.435 118.715 20.665 ;
        RECT 119.635 20.435 120.875 20.665 ;
        RECT 117.475 19.740 117.735 20.435 ;
        RECT 111.860 19.140 112.870 19.310 ;
        RECT 111.860 17.180 112.030 19.140 ;
        RECT 112.190 17.625 112.450 18.760 ;
        RECT 112.640 17.830 112.870 19.140 ;
        RECT 113.415 19.080 113.675 19.400 ;
        RECT 114.005 19.080 114.265 19.400 ;
        RECT 114.795 19.080 115.055 19.400 ;
        RECT 113.430 17.830 113.660 19.080 ;
        RECT 114.020 17.830 114.250 19.080 ;
        RECT 114.810 17.830 115.040 19.080 ;
        RECT 115.280 17.625 115.540 18.130 ;
        RECT 112.190 17.395 113.380 17.625 ;
        RECT 114.300 17.395 115.540 17.625 ;
        RECT 115.965 17.180 116.320 19.370 ;
        RECT 111.365 16.905 112.030 17.180 ;
        RECT 115.650 16.905 116.320 17.180 ;
        RECT 111.365 14.800 111.720 16.905 ;
        RECT 112.140 16.480 113.380 16.710 ;
        RECT 114.300 16.480 115.490 16.710 ;
        RECT 112.140 16.055 112.400 16.480 ;
        RECT 112.640 15.040 112.870 16.275 ;
        RECT 113.430 15.040 113.660 16.275 ;
        RECT 114.020 15.040 114.250 16.275 ;
        RECT 104.620 13.670 104.880 14.460 ;
        RECT 101.480 13.440 102.720 13.670 ;
        RECT 103.640 13.440 104.880 13.670 ;
        RECT 106.815 13.670 107.075 14.550 ;
        RECT 107.315 13.830 107.545 14.720 ;
        RECT 108.105 13.830 108.335 14.720 ;
        RECT 108.695 13.830 108.925 14.720 ;
        RECT 109.485 13.830 109.715 14.795 ;
        RECT 112.625 14.720 112.885 15.040 ;
        RECT 113.415 14.720 113.675 15.040 ;
        RECT 114.005 14.720 114.265 15.040 ;
        RECT 114.810 14.965 115.040 16.275 ;
        RECT 115.230 15.405 115.490 16.480 ;
        RECT 115.650 14.965 115.820 16.905 ;
        RECT 114.810 14.795 115.820 14.965 ;
        RECT 115.965 14.795 116.320 16.905 ;
        RECT 116.700 17.180 117.055 19.375 ;
        RECT 117.975 19.310 118.205 20.275 ;
        RECT 118.765 19.400 118.995 20.275 ;
        RECT 119.355 19.400 119.585 20.275 ;
        RECT 120.145 19.400 120.375 20.275 ;
        RECT 120.615 19.645 120.875 20.435 ;
        RECT 117.195 19.140 118.205 19.310 ;
        RECT 117.195 17.180 117.365 19.140 ;
        RECT 117.525 17.625 117.785 18.760 ;
        RECT 117.975 17.830 118.205 19.140 ;
        RECT 118.750 19.080 119.010 19.400 ;
        RECT 119.340 19.080 119.600 19.400 ;
        RECT 120.130 19.080 120.390 19.400 ;
        RECT 118.765 17.830 118.995 19.080 ;
        RECT 119.355 17.830 119.585 19.080 ;
        RECT 120.145 17.830 120.375 19.080 ;
        RECT 120.615 17.625 120.875 18.130 ;
        RECT 117.525 17.395 118.715 17.625 ;
        RECT 119.635 17.395 120.875 17.625 ;
        RECT 121.300 17.180 121.655 19.370 ;
        RECT 116.700 16.905 117.365 17.180 ;
        RECT 120.985 16.905 121.655 17.180 ;
        RECT 116.700 14.800 117.055 16.905 ;
        RECT 117.475 16.480 118.715 16.710 ;
        RECT 119.635 16.480 120.825 16.710 ;
        RECT 117.475 16.055 117.735 16.480 ;
        RECT 117.975 15.040 118.205 16.275 ;
        RECT 118.765 15.040 118.995 16.275 ;
        RECT 119.355 15.040 119.585 16.275 ;
        RECT 109.955 13.670 110.215 14.460 ;
        RECT 106.815 13.440 108.055 13.670 ;
        RECT 108.975 13.440 110.215 13.670 ;
        RECT 112.140 13.670 112.400 14.550 ;
        RECT 112.640 13.830 112.870 14.720 ;
        RECT 113.430 13.830 113.660 14.720 ;
        RECT 114.020 13.830 114.250 14.720 ;
        RECT 114.810 13.830 115.040 14.795 ;
        RECT 117.960 14.720 118.220 15.040 ;
        RECT 118.750 14.720 119.010 15.040 ;
        RECT 119.340 14.720 119.600 15.040 ;
        RECT 120.145 14.965 120.375 16.275 ;
        RECT 120.565 15.405 120.825 16.480 ;
        RECT 120.985 14.965 121.155 16.905 ;
        RECT 120.145 14.795 121.155 14.965 ;
        RECT 121.300 14.795 121.655 16.905 ;
        RECT 122.025 17.180 122.380 19.390 ;
        RECT 123.300 19.310 123.530 20.275 ;
        RECT 124.090 19.400 124.320 20.275 ;
        RECT 124.680 19.400 124.910 20.275 ;
        RECT 125.470 19.400 125.700 20.275 ;
        RECT 122.520 19.140 123.530 19.310 ;
        RECT 122.520 17.180 122.690 19.140 ;
        RECT 123.300 17.830 123.530 19.140 ;
        RECT 124.075 19.080 124.335 19.400 ;
        RECT 124.665 19.080 124.925 19.400 ;
        RECT 125.455 19.080 125.715 19.400 ;
        RECT 124.090 17.830 124.320 19.080 ;
        RECT 124.680 17.830 124.910 19.080 ;
        RECT 125.470 17.830 125.700 19.080 ;
        RECT 126.625 17.180 126.980 19.390 ;
        RECT 122.025 16.905 122.690 17.180 ;
        RECT 126.310 16.905 126.980 17.180 ;
        RECT 122.025 14.815 122.380 16.905 ;
        RECT 123.300 15.040 123.530 16.275 ;
        RECT 124.090 15.040 124.320 16.275 ;
        RECT 124.680 15.040 124.910 16.275 ;
        RECT 115.280 13.670 115.540 14.460 ;
        RECT 112.140 13.440 113.380 13.670 ;
        RECT 114.300 13.440 115.540 13.670 ;
        RECT 117.475 13.670 117.735 14.550 ;
        RECT 117.975 13.830 118.205 14.720 ;
        RECT 118.765 13.830 118.995 14.720 ;
        RECT 119.355 13.830 119.585 14.720 ;
        RECT 120.145 13.830 120.375 14.795 ;
        RECT 123.285 14.720 123.545 15.040 ;
        RECT 124.075 14.720 124.335 15.040 ;
        RECT 124.665 14.720 124.925 15.040 ;
        RECT 125.470 14.965 125.700 16.275 ;
        RECT 126.310 14.965 126.480 16.905 ;
        RECT 125.470 14.795 126.480 14.965 ;
        RECT 126.625 14.815 126.980 16.905 ;
        RECT 120.615 13.670 120.875 14.460 ;
        RECT 123.300 13.830 123.530 14.720 ;
        RECT 124.090 13.830 124.320 14.720 ;
        RECT 124.680 13.830 124.910 14.720 ;
        RECT 125.470 13.830 125.700 14.795 ;
        RECT 117.475 13.440 118.715 13.670 ;
        RECT 119.635 13.440 120.875 13.670 ;
        RECT 37.520 12.900 38.760 13.130 ;
        RECT 39.680 12.900 40.920 13.130 ;
        RECT 10.500 11.770 10.820 12.255 ;
        RECT 16.115 11.880 27.620 12.115 ;
        RECT 10.500 11.440 11.960 11.770 ;
        RECT 10.500 11.220 10.820 11.440 ;
        RECT 12.400 10.695 12.720 11.685 ;
        RECT 14.585 11.440 16.005 11.765 ;
        RECT 19.990 11.310 27.620 11.880 ;
        RECT 16.115 11.075 27.620 11.310 ;
        RECT 12.425 10.680 12.715 10.695 ;
        RECT 31.420 10.230 31.775 11.855 ;
        RECT 32.695 11.775 32.925 12.740 ;
        RECT 33.485 11.865 33.715 12.740 ;
        RECT 34.075 11.865 34.305 12.740 ;
        RECT 34.865 11.865 35.095 12.740 ;
        RECT 37.520 12.205 37.780 12.900 ;
        RECT 38.810 11.865 39.040 12.740 ;
        RECT 39.400 11.865 39.630 12.740 ;
        RECT 40.190 11.865 40.420 12.740 ;
        RECT 40.660 12.110 40.920 12.900 ;
        RECT 42.855 12.900 44.095 13.130 ;
        RECT 45.015 12.900 46.255 13.130 ;
        RECT 42.855 12.205 43.115 12.900 ;
        RECT 31.240 9.645 31.775 10.230 ;
        RECT 31.915 11.605 32.925 11.775 ;
        RECT 31.915 9.645 32.085 11.605 ;
        RECT 32.695 10.295 32.925 11.605 ;
        RECT 33.470 11.545 33.730 11.865 ;
        RECT 34.060 11.545 34.320 11.865 ;
        RECT 34.850 11.545 35.110 11.865 ;
        RECT 38.795 11.545 39.055 11.865 ;
        RECT 39.385 11.545 39.645 11.865 ;
        RECT 40.175 11.545 40.435 11.865 ;
        RECT 33.485 10.295 33.715 11.545 ;
        RECT 34.075 10.295 34.305 11.545 ;
        RECT 34.865 10.295 35.095 11.545 ;
        RECT 37.570 10.090 37.830 11.225 ;
        RECT 38.810 10.295 39.040 11.545 ;
        RECT 39.400 10.295 39.630 11.545 ;
        RECT 40.190 10.295 40.420 11.545 ;
        RECT 40.660 10.090 40.920 10.595 ;
        RECT 37.570 9.860 38.760 10.090 ;
        RECT 39.680 9.860 40.920 10.090 ;
        RECT 41.345 10.230 41.700 11.835 ;
        RECT 42.080 10.230 42.435 11.840 ;
        RECT 43.355 11.775 43.585 12.740 ;
        RECT 44.145 11.865 44.375 12.740 ;
        RECT 44.735 11.865 44.965 12.740 ;
        RECT 45.525 11.865 45.755 12.740 ;
        RECT 45.995 12.110 46.255 12.900 ;
        RECT 48.180 12.900 49.420 13.130 ;
        RECT 50.340 12.900 51.580 13.130 ;
        RECT 48.180 12.205 48.440 12.900 ;
        RECT 41.345 9.645 42.435 10.230 ;
        RECT 42.575 11.605 43.585 11.775 ;
        RECT 42.575 9.645 42.745 11.605 ;
        RECT 42.905 10.090 43.165 11.225 ;
        RECT 43.355 10.295 43.585 11.605 ;
        RECT 44.130 11.545 44.390 11.865 ;
        RECT 44.720 11.545 44.980 11.865 ;
        RECT 45.510 11.545 45.770 11.865 ;
        RECT 44.145 10.295 44.375 11.545 ;
        RECT 44.735 10.295 44.965 11.545 ;
        RECT 45.525 10.295 45.755 11.545 ;
        RECT 45.995 10.090 46.255 10.595 ;
        RECT 42.905 9.860 44.095 10.090 ;
        RECT 45.015 9.860 46.255 10.090 ;
        RECT 46.680 10.235 47.035 11.835 ;
        RECT 47.405 10.235 47.760 11.840 ;
        RECT 48.680 11.775 48.910 12.740 ;
        RECT 49.470 11.865 49.700 12.740 ;
        RECT 50.060 11.865 50.290 12.740 ;
        RECT 50.850 11.865 51.080 12.740 ;
        RECT 51.320 12.110 51.580 12.900 ;
        RECT 53.515 12.900 54.755 13.130 ;
        RECT 55.675 12.900 56.915 13.130 ;
        RECT 53.515 12.205 53.775 12.900 ;
        RECT 46.680 9.650 47.760 10.235 ;
        RECT 46.680 9.645 47.035 9.650 ;
        RECT 31.420 9.370 32.085 9.645 ;
        RECT 41.030 9.370 41.700 9.645 ;
        RECT 15.985 8.690 22.260 8.695 ;
        RECT 28.045 8.690 28.305 8.695 ;
        RECT 10.510 7.175 10.810 8.625 ;
        RECT 15.985 8.460 28.345 8.690 ;
        RECT 11.745 8.075 13.345 8.365 ;
        RECT 14.165 8.075 20.945 8.310 ;
        RECT 16.040 7.890 17.645 7.920 ;
        RECT 21.425 7.890 28.345 8.460 ;
        RECT 15.985 7.655 28.345 7.890 ;
        RECT 16.040 7.630 17.645 7.655 ;
        RECT 31.420 7.280 31.775 9.370 ;
        RECT 32.695 7.505 32.925 8.740 ;
        RECT 33.485 7.505 33.715 8.740 ;
        RECT 34.075 7.505 34.305 8.740 ;
        RECT 38.020 7.505 38.250 8.740 ;
        RECT 38.810 7.505 39.040 8.740 ;
        RECT 39.400 7.505 39.630 8.740 ;
        RECT 31.460 4.320 31.710 7.280 ;
        RECT 32.680 7.185 32.940 7.505 ;
        RECT 33.470 7.185 33.730 7.505 ;
        RECT 34.060 7.185 34.320 7.505 ;
        RECT 38.005 7.185 38.265 7.505 ;
        RECT 38.795 7.185 39.055 7.505 ;
        RECT 39.385 7.185 39.645 7.505 ;
        RECT 40.190 7.430 40.420 8.740 ;
        RECT 41.030 7.430 41.200 9.370 ;
        RECT 40.190 7.260 41.200 7.430 ;
        RECT 41.345 7.260 41.700 9.370 ;
        RECT 42.080 9.370 42.745 9.645 ;
        RECT 46.365 9.370 47.035 9.645 ;
        RECT 42.080 7.265 42.435 9.370 ;
        RECT 43.355 7.505 43.585 8.740 ;
        RECT 44.145 7.505 44.375 8.740 ;
        RECT 44.735 7.505 44.965 8.740 ;
        RECT 32.695 6.295 32.925 7.185 ;
        RECT 33.485 6.295 33.715 7.185 ;
        RECT 34.075 6.295 34.305 7.185 ;
        RECT 38.020 6.295 38.250 7.185 ;
        RECT 38.810 6.295 39.040 7.185 ;
        RECT 39.400 6.295 39.630 7.185 ;
        RECT 40.190 6.295 40.420 7.260 ;
        RECT 43.340 7.185 43.600 7.505 ;
        RECT 44.130 7.185 44.390 7.505 ;
        RECT 44.720 7.185 44.980 7.505 ;
        RECT 45.525 7.430 45.755 8.740 ;
        RECT 46.365 7.430 46.535 9.370 ;
        RECT 45.525 7.260 46.535 7.430 ;
        RECT 46.680 7.260 47.035 9.370 ;
        RECT 47.405 9.645 47.760 9.650 ;
        RECT 47.900 11.605 48.910 11.775 ;
        RECT 47.900 9.645 48.070 11.605 ;
        RECT 48.230 10.090 48.490 11.225 ;
        RECT 48.680 10.295 48.910 11.605 ;
        RECT 49.455 11.545 49.715 11.865 ;
        RECT 50.045 11.545 50.305 11.865 ;
        RECT 50.835 11.545 51.095 11.865 ;
        RECT 49.470 10.295 49.700 11.545 ;
        RECT 50.060 10.295 50.290 11.545 ;
        RECT 50.850 10.295 51.080 11.545 ;
        RECT 51.320 10.090 51.580 10.595 ;
        RECT 48.230 9.860 49.420 10.090 ;
        RECT 50.340 9.860 51.580 10.090 ;
        RECT 52.005 10.230 52.360 11.835 ;
        RECT 52.740 10.230 53.095 11.840 ;
        RECT 54.015 11.775 54.245 12.740 ;
        RECT 54.805 11.865 55.035 12.740 ;
        RECT 55.395 11.865 55.625 12.740 ;
        RECT 56.185 11.865 56.415 12.740 ;
        RECT 56.655 12.110 56.915 12.900 ;
        RECT 58.840 12.900 60.080 13.130 ;
        RECT 61.000 12.900 62.240 13.130 ;
        RECT 58.840 12.205 59.100 12.900 ;
        RECT 52.005 9.645 53.095 10.230 ;
        RECT 53.235 11.605 54.245 11.775 ;
        RECT 53.235 9.645 53.405 11.605 ;
        RECT 53.565 10.090 53.825 11.225 ;
        RECT 54.015 10.295 54.245 11.605 ;
        RECT 54.790 11.545 55.050 11.865 ;
        RECT 55.380 11.545 55.640 11.865 ;
        RECT 56.170 11.545 56.430 11.865 ;
        RECT 54.805 10.295 55.035 11.545 ;
        RECT 55.395 10.295 55.625 11.545 ;
        RECT 56.185 10.295 56.415 11.545 ;
        RECT 56.655 10.090 56.915 10.595 ;
        RECT 53.565 9.860 54.755 10.090 ;
        RECT 55.675 9.860 56.915 10.090 ;
        RECT 57.340 10.235 57.695 11.835 ;
        RECT 58.065 10.235 58.420 11.840 ;
        RECT 59.340 11.775 59.570 12.740 ;
        RECT 60.130 11.865 60.360 12.740 ;
        RECT 60.720 11.865 60.950 12.740 ;
        RECT 61.510 11.865 61.740 12.740 ;
        RECT 61.980 12.110 62.240 12.900 ;
        RECT 64.175 12.900 65.415 13.130 ;
        RECT 66.335 12.900 67.575 13.130 ;
        RECT 64.175 12.205 64.435 12.900 ;
        RECT 57.340 9.650 58.420 10.235 ;
        RECT 57.340 9.645 57.695 9.650 ;
        RECT 47.405 9.370 48.070 9.645 ;
        RECT 51.690 9.370 52.360 9.645 ;
        RECT 47.405 7.265 47.760 9.370 ;
        RECT 48.680 7.505 48.910 8.740 ;
        RECT 49.470 7.505 49.700 8.740 ;
        RECT 50.060 7.505 50.290 8.740 ;
        RECT 43.355 6.295 43.585 7.185 ;
        RECT 44.145 6.295 44.375 7.185 ;
        RECT 44.735 6.295 44.965 7.185 ;
        RECT 45.525 6.295 45.755 7.260 ;
        RECT 48.665 7.185 48.925 7.505 ;
        RECT 49.455 7.185 49.715 7.505 ;
        RECT 50.045 7.185 50.305 7.505 ;
        RECT 50.850 7.430 51.080 8.740 ;
        RECT 51.690 7.430 51.860 9.370 ;
        RECT 50.850 7.260 51.860 7.430 ;
        RECT 52.005 7.260 52.360 9.370 ;
        RECT 52.740 9.370 53.405 9.645 ;
        RECT 57.025 9.370 57.695 9.645 ;
        RECT 52.740 7.265 53.095 9.370 ;
        RECT 54.015 7.505 54.245 8.740 ;
        RECT 54.805 7.505 55.035 8.740 ;
        RECT 55.395 7.505 55.625 8.740 ;
        RECT 48.680 6.295 48.910 7.185 ;
        RECT 49.470 6.295 49.700 7.185 ;
        RECT 50.060 6.295 50.290 7.185 ;
        RECT 50.850 6.295 51.080 7.260 ;
        RECT 54.000 7.185 54.260 7.505 ;
        RECT 54.790 7.185 55.050 7.505 ;
        RECT 55.380 7.185 55.640 7.505 ;
        RECT 56.185 7.430 56.415 8.740 ;
        RECT 57.025 7.430 57.195 9.370 ;
        RECT 56.185 7.260 57.195 7.430 ;
        RECT 57.340 7.260 57.695 9.370 ;
        RECT 58.065 9.645 58.420 9.650 ;
        RECT 58.560 11.605 59.570 11.775 ;
        RECT 58.560 9.645 58.730 11.605 ;
        RECT 58.890 10.090 59.150 11.225 ;
        RECT 59.340 10.295 59.570 11.605 ;
        RECT 60.115 11.545 60.375 11.865 ;
        RECT 60.705 11.545 60.965 11.865 ;
        RECT 61.495 11.545 61.755 11.865 ;
        RECT 60.130 10.295 60.360 11.545 ;
        RECT 60.720 10.295 60.950 11.545 ;
        RECT 61.510 10.295 61.740 11.545 ;
        RECT 61.980 10.090 62.240 10.595 ;
        RECT 58.890 9.860 60.080 10.090 ;
        RECT 61.000 9.860 62.240 10.090 ;
        RECT 62.665 10.230 63.020 11.835 ;
        RECT 63.400 10.230 63.755 11.840 ;
        RECT 64.675 11.775 64.905 12.740 ;
        RECT 65.465 11.865 65.695 12.740 ;
        RECT 66.055 11.865 66.285 12.740 ;
        RECT 66.845 11.865 67.075 12.740 ;
        RECT 67.315 12.110 67.575 12.900 ;
        RECT 69.500 12.900 70.740 13.130 ;
        RECT 71.660 12.900 72.900 13.130 ;
        RECT 69.500 12.205 69.760 12.900 ;
        RECT 62.665 9.645 63.755 10.230 ;
        RECT 63.895 11.605 64.905 11.775 ;
        RECT 63.895 9.645 64.065 11.605 ;
        RECT 64.225 10.090 64.485 11.225 ;
        RECT 64.675 10.295 64.905 11.605 ;
        RECT 65.450 11.545 65.710 11.865 ;
        RECT 66.040 11.545 66.300 11.865 ;
        RECT 66.830 11.545 67.090 11.865 ;
        RECT 65.465 10.295 65.695 11.545 ;
        RECT 66.055 10.295 66.285 11.545 ;
        RECT 66.845 10.295 67.075 11.545 ;
        RECT 67.315 10.090 67.575 10.595 ;
        RECT 64.225 9.860 65.415 10.090 ;
        RECT 66.335 9.860 67.575 10.090 ;
        RECT 68.000 10.235 68.355 11.835 ;
        RECT 68.725 10.235 69.080 11.840 ;
        RECT 70.000 11.775 70.230 12.740 ;
        RECT 70.790 11.865 71.020 12.740 ;
        RECT 71.380 11.865 71.610 12.740 ;
        RECT 72.170 11.865 72.400 12.740 ;
        RECT 72.640 12.110 72.900 12.900 ;
        RECT 74.835 12.900 76.075 13.130 ;
        RECT 76.995 12.900 78.235 13.130 ;
        RECT 74.835 12.205 75.095 12.900 ;
        RECT 68.000 9.650 69.080 10.235 ;
        RECT 68.000 9.645 68.355 9.650 ;
        RECT 58.065 9.370 58.730 9.645 ;
        RECT 62.350 9.370 63.020 9.645 ;
        RECT 58.065 7.265 58.420 9.370 ;
        RECT 59.340 7.505 59.570 8.740 ;
        RECT 60.130 7.505 60.360 8.740 ;
        RECT 60.720 7.505 60.950 8.740 ;
        RECT 54.015 6.295 54.245 7.185 ;
        RECT 54.805 6.295 55.035 7.185 ;
        RECT 55.395 6.295 55.625 7.185 ;
        RECT 56.185 6.295 56.415 7.260 ;
        RECT 59.325 7.185 59.585 7.505 ;
        RECT 60.115 7.185 60.375 7.505 ;
        RECT 60.705 7.185 60.965 7.505 ;
        RECT 61.510 7.430 61.740 8.740 ;
        RECT 62.350 7.430 62.520 9.370 ;
        RECT 61.510 7.260 62.520 7.430 ;
        RECT 62.665 7.260 63.020 9.370 ;
        RECT 63.400 9.370 64.065 9.645 ;
        RECT 67.685 9.370 68.355 9.645 ;
        RECT 63.400 7.265 63.755 9.370 ;
        RECT 64.675 7.505 64.905 8.740 ;
        RECT 65.465 7.505 65.695 8.740 ;
        RECT 66.055 7.505 66.285 8.740 ;
        RECT 59.340 6.295 59.570 7.185 ;
        RECT 60.130 6.295 60.360 7.185 ;
        RECT 60.720 6.295 60.950 7.185 ;
        RECT 61.510 6.295 61.740 7.260 ;
        RECT 64.660 7.185 64.920 7.505 ;
        RECT 65.450 7.185 65.710 7.505 ;
        RECT 66.040 7.185 66.300 7.505 ;
        RECT 66.845 7.430 67.075 8.740 ;
        RECT 67.685 7.430 67.855 9.370 ;
        RECT 66.845 7.260 67.855 7.430 ;
        RECT 68.000 7.260 68.355 9.370 ;
        RECT 68.725 9.645 69.080 9.650 ;
        RECT 69.220 11.605 70.230 11.775 ;
        RECT 69.220 9.645 69.390 11.605 ;
        RECT 69.550 10.090 69.810 11.225 ;
        RECT 70.000 10.295 70.230 11.605 ;
        RECT 70.775 11.545 71.035 11.865 ;
        RECT 71.365 11.545 71.625 11.865 ;
        RECT 72.155 11.545 72.415 11.865 ;
        RECT 70.790 10.295 71.020 11.545 ;
        RECT 71.380 10.295 71.610 11.545 ;
        RECT 72.170 10.295 72.400 11.545 ;
        RECT 72.640 10.090 72.900 10.595 ;
        RECT 69.550 9.860 70.740 10.090 ;
        RECT 71.660 9.860 72.900 10.090 ;
        RECT 73.325 10.230 73.680 11.835 ;
        RECT 74.060 10.230 74.415 11.840 ;
        RECT 75.335 11.775 75.565 12.740 ;
        RECT 76.125 11.865 76.355 12.740 ;
        RECT 76.715 11.865 76.945 12.740 ;
        RECT 77.505 11.865 77.735 12.740 ;
        RECT 77.975 12.110 78.235 12.900 ;
        RECT 80.160 12.900 81.400 13.130 ;
        RECT 82.320 12.900 83.560 13.130 ;
        RECT 80.160 12.205 80.420 12.900 ;
        RECT 73.325 9.645 74.415 10.230 ;
        RECT 74.555 11.605 75.565 11.775 ;
        RECT 74.555 9.645 74.725 11.605 ;
        RECT 74.885 10.090 75.145 11.225 ;
        RECT 75.335 10.295 75.565 11.605 ;
        RECT 76.110 11.545 76.370 11.865 ;
        RECT 76.700 11.545 76.960 11.865 ;
        RECT 77.490 11.545 77.750 11.865 ;
        RECT 76.125 10.295 76.355 11.545 ;
        RECT 76.715 10.295 76.945 11.545 ;
        RECT 77.505 10.295 77.735 11.545 ;
        RECT 77.975 10.090 78.235 10.595 ;
        RECT 74.885 9.860 76.075 10.090 ;
        RECT 76.995 9.860 78.235 10.090 ;
        RECT 78.660 10.235 79.015 11.835 ;
        RECT 79.385 10.235 79.740 11.840 ;
        RECT 80.660 11.775 80.890 12.740 ;
        RECT 81.450 11.865 81.680 12.740 ;
        RECT 82.040 11.865 82.270 12.740 ;
        RECT 82.830 11.865 83.060 12.740 ;
        RECT 83.300 12.110 83.560 12.900 ;
        RECT 85.495 12.900 86.735 13.130 ;
        RECT 87.655 12.900 88.895 13.130 ;
        RECT 85.495 12.205 85.755 12.900 ;
        RECT 78.660 9.650 79.740 10.235 ;
        RECT 78.660 9.645 79.015 9.650 ;
        RECT 68.725 9.370 69.390 9.645 ;
        RECT 73.010 9.370 73.680 9.645 ;
        RECT 68.725 7.265 69.080 9.370 ;
        RECT 70.000 7.505 70.230 8.740 ;
        RECT 70.790 7.505 71.020 8.740 ;
        RECT 71.380 7.505 71.610 8.740 ;
        RECT 64.675 6.295 64.905 7.185 ;
        RECT 65.465 6.295 65.695 7.185 ;
        RECT 66.055 6.295 66.285 7.185 ;
        RECT 66.845 6.295 67.075 7.260 ;
        RECT 69.985 7.185 70.245 7.505 ;
        RECT 70.775 7.185 71.035 7.505 ;
        RECT 71.365 7.185 71.625 7.505 ;
        RECT 72.170 7.430 72.400 8.740 ;
        RECT 73.010 7.430 73.180 9.370 ;
        RECT 72.170 7.260 73.180 7.430 ;
        RECT 73.325 7.260 73.680 9.370 ;
        RECT 74.060 9.370 74.725 9.645 ;
        RECT 78.345 9.370 79.015 9.645 ;
        RECT 74.060 7.265 74.415 9.370 ;
        RECT 75.335 7.505 75.565 8.740 ;
        RECT 76.125 7.505 76.355 8.740 ;
        RECT 76.715 7.505 76.945 8.740 ;
        RECT 70.000 6.295 70.230 7.185 ;
        RECT 70.790 6.295 71.020 7.185 ;
        RECT 71.380 6.295 71.610 7.185 ;
        RECT 72.170 6.295 72.400 7.260 ;
        RECT 75.320 7.185 75.580 7.505 ;
        RECT 76.110 7.185 76.370 7.505 ;
        RECT 76.700 7.185 76.960 7.505 ;
        RECT 77.505 7.430 77.735 8.740 ;
        RECT 78.345 7.430 78.515 9.370 ;
        RECT 77.505 7.260 78.515 7.430 ;
        RECT 78.660 7.260 79.015 9.370 ;
        RECT 79.385 9.645 79.740 9.650 ;
        RECT 79.880 11.605 80.890 11.775 ;
        RECT 79.880 9.645 80.050 11.605 ;
        RECT 80.210 10.090 80.470 11.225 ;
        RECT 80.660 10.295 80.890 11.605 ;
        RECT 81.435 11.545 81.695 11.865 ;
        RECT 82.025 11.545 82.285 11.865 ;
        RECT 82.815 11.545 83.075 11.865 ;
        RECT 81.450 10.295 81.680 11.545 ;
        RECT 82.040 10.295 82.270 11.545 ;
        RECT 82.830 10.295 83.060 11.545 ;
        RECT 83.300 10.090 83.560 10.595 ;
        RECT 80.210 9.860 81.400 10.090 ;
        RECT 82.320 9.860 83.560 10.090 ;
        RECT 83.985 10.230 84.340 11.835 ;
        RECT 84.720 10.230 85.075 11.840 ;
        RECT 85.995 11.775 86.225 12.740 ;
        RECT 86.785 11.865 87.015 12.740 ;
        RECT 87.375 11.865 87.605 12.740 ;
        RECT 88.165 11.865 88.395 12.740 ;
        RECT 88.635 12.110 88.895 12.900 ;
        RECT 90.820 12.900 92.060 13.130 ;
        RECT 92.980 12.900 94.220 13.130 ;
        RECT 90.820 12.205 91.080 12.900 ;
        RECT 83.985 9.645 85.075 10.230 ;
        RECT 85.215 11.605 86.225 11.775 ;
        RECT 85.215 9.645 85.385 11.605 ;
        RECT 85.545 10.090 85.805 11.225 ;
        RECT 85.995 10.295 86.225 11.605 ;
        RECT 86.770 11.545 87.030 11.865 ;
        RECT 87.360 11.545 87.620 11.865 ;
        RECT 88.150 11.545 88.410 11.865 ;
        RECT 86.785 10.295 87.015 11.545 ;
        RECT 87.375 10.295 87.605 11.545 ;
        RECT 88.165 10.295 88.395 11.545 ;
        RECT 88.635 10.090 88.895 10.595 ;
        RECT 85.545 9.860 86.735 10.090 ;
        RECT 87.655 9.860 88.895 10.090 ;
        RECT 89.320 10.235 89.675 11.835 ;
        RECT 90.045 10.235 90.400 11.840 ;
        RECT 91.320 11.775 91.550 12.740 ;
        RECT 92.110 11.865 92.340 12.740 ;
        RECT 92.700 11.865 92.930 12.740 ;
        RECT 93.490 11.865 93.720 12.740 ;
        RECT 93.960 12.110 94.220 12.900 ;
        RECT 96.155 12.900 97.395 13.130 ;
        RECT 98.315 12.900 99.555 13.130 ;
        RECT 96.155 12.205 96.415 12.900 ;
        RECT 89.320 9.650 90.400 10.235 ;
        RECT 89.320 9.645 89.675 9.650 ;
        RECT 79.385 9.370 80.050 9.645 ;
        RECT 83.670 9.370 84.340 9.645 ;
        RECT 79.385 7.265 79.740 9.370 ;
        RECT 80.660 7.505 80.890 8.740 ;
        RECT 81.450 7.505 81.680 8.740 ;
        RECT 82.040 7.505 82.270 8.740 ;
        RECT 75.335 6.295 75.565 7.185 ;
        RECT 76.125 6.295 76.355 7.185 ;
        RECT 76.715 6.295 76.945 7.185 ;
        RECT 77.505 6.295 77.735 7.260 ;
        RECT 80.645 7.185 80.905 7.505 ;
        RECT 81.435 7.185 81.695 7.505 ;
        RECT 82.025 7.185 82.285 7.505 ;
        RECT 82.830 7.430 83.060 8.740 ;
        RECT 83.670 7.430 83.840 9.370 ;
        RECT 82.830 7.260 83.840 7.430 ;
        RECT 83.985 7.260 84.340 9.370 ;
        RECT 84.720 9.370 85.385 9.645 ;
        RECT 89.005 9.370 89.675 9.645 ;
        RECT 84.720 7.265 85.075 9.370 ;
        RECT 85.995 7.505 86.225 8.740 ;
        RECT 86.785 7.505 87.015 8.740 ;
        RECT 87.375 7.505 87.605 8.740 ;
        RECT 80.660 6.295 80.890 7.185 ;
        RECT 81.450 6.295 81.680 7.185 ;
        RECT 82.040 6.295 82.270 7.185 ;
        RECT 82.830 6.295 83.060 7.260 ;
        RECT 85.980 7.185 86.240 7.505 ;
        RECT 86.770 7.185 87.030 7.505 ;
        RECT 87.360 7.185 87.620 7.505 ;
        RECT 88.165 7.430 88.395 8.740 ;
        RECT 89.005 7.430 89.175 9.370 ;
        RECT 88.165 7.260 89.175 7.430 ;
        RECT 89.320 7.260 89.675 9.370 ;
        RECT 90.045 9.645 90.400 9.650 ;
        RECT 90.540 11.605 91.550 11.775 ;
        RECT 90.540 9.645 90.710 11.605 ;
        RECT 90.870 10.090 91.130 11.225 ;
        RECT 91.320 10.295 91.550 11.605 ;
        RECT 92.095 11.545 92.355 11.865 ;
        RECT 92.685 11.545 92.945 11.865 ;
        RECT 93.475 11.545 93.735 11.865 ;
        RECT 92.110 10.295 92.340 11.545 ;
        RECT 92.700 10.295 92.930 11.545 ;
        RECT 93.490 10.295 93.720 11.545 ;
        RECT 93.960 10.090 94.220 10.595 ;
        RECT 90.870 9.860 92.060 10.090 ;
        RECT 92.980 9.860 94.220 10.090 ;
        RECT 94.645 10.230 95.000 11.835 ;
        RECT 95.380 10.230 95.735 11.840 ;
        RECT 96.655 11.775 96.885 12.740 ;
        RECT 97.445 11.865 97.675 12.740 ;
        RECT 98.035 11.865 98.265 12.740 ;
        RECT 98.825 11.865 99.055 12.740 ;
        RECT 99.295 12.110 99.555 12.900 ;
        RECT 101.480 12.900 102.720 13.130 ;
        RECT 103.640 12.900 104.880 13.130 ;
        RECT 101.480 12.205 101.740 12.900 ;
        RECT 94.645 9.645 95.735 10.230 ;
        RECT 95.875 11.605 96.885 11.775 ;
        RECT 95.875 9.645 96.045 11.605 ;
        RECT 96.205 10.090 96.465 11.225 ;
        RECT 96.655 10.295 96.885 11.605 ;
        RECT 97.430 11.545 97.690 11.865 ;
        RECT 98.020 11.545 98.280 11.865 ;
        RECT 98.810 11.545 99.070 11.865 ;
        RECT 97.445 10.295 97.675 11.545 ;
        RECT 98.035 10.295 98.265 11.545 ;
        RECT 98.825 10.295 99.055 11.545 ;
        RECT 99.295 10.090 99.555 10.595 ;
        RECT 96.205 9.860 97.395 10.090 ;
        RECT 98.315 9.860 99.555 10.090 ;
        RECT 99.980 10.235 100.335 11.835 ;
        RECT 100.705 10.235 101.060 11.840 ;
        RECT 101.980 11.775 102.210 12.740 ;
        RECT 102.770 11.865 103.000 12.740 ;
        RECT 103.360 11.865 103.590 12.740 ;
        RECT 104.150 11.865 104.380 12.740 ;
        RECT 104.620 12.110 104.880 12.900 ;
        RECT 106.815 12.900 108.055 13.130 ;
        RECT 108.975 12.900 110.215 13.130 ;
        RECT 106.815 12.205 107.075 12.900 ;
        RECT 99.980 9.650 101.060 10.235 ;
        RECT 99.980 9.645 100.335 9.650 ;
        RECT 90.045 9.370 90.710 9.645 ;
        RECT 94.330 9.370 95.000 9.645 ;
        RECT 90.045 7.265 90.400 9.370 ;
        RECT 91.320 7.505 91.550 8.740 ;
        RECT 92.110 7.505 92.340 8.740 ;
        RECT 92.700 7.505 92.930 8.740 ;
        RECT 85.995 6.295 86.225 7.185 ;
        RECT 86.785 6.295 87.015 7.185 ;
        RECT 87.375 6.295 87.605 7.185 ;
        RECT 88.165 6.295 88.395 7.260 ;
        RECT 91.305 7.185 91.565 7.505 ;
        RECT 92.095 7.185 92.355 7.505 ;
        RECT 92.685 7.185 92.945 7.505 ;
        RECT 93.490 7.430 93.720 8.740 ;
        RECT 94.330 7.430 94.500 9.370 ;
        RECT 93.490 7.260 94.500 7.430 ;
        RECT 94.645 7.260 95.000 9.370 ;
        RECT 95.380 9.370 96.045 9.645 ;
        RECT 99.665 9.370 100.335 9.645 ;
        RECT 95.380 7.265 95.735 9.370 ;
        RECT 96.655 7.505 96.885 8.740 ;
        RECT 97.445 7.505 97.675 8.740 ;
        RECT 98.035 7.505 98.265 8.740 ;
        RECT 91.320 6.295 91.550 7.185 ;
        RECT 92.110 6.295 92.340 7.185 ;
        RECT 92.700 6.295 92.930 7.185 ;
        RECT 93.490 6.295 93.720 7.260 ;
        RECT 96.640 7.185 96.900 7.505 ;
        RECT 97.430 7.185 97.690 7.505 ;
        RECT 98.020 7.185 98.280 7.505 ;
        RECT 98.825 7.430 99.055 8.740 ;
        RECT 99.665 7.430 99.835 9.370 ;
        RECT 98.825 7.260 99.835 7.430 ;
        RECT 99.980 7.260 100.335 9.370 ;
        RECT 100.705 9.645 101.060 9.650 ;
        RECT 101.200 11.605 102.210 11.775 ;
        RECT 101.200 9.645 101.370 11.605 ;
        RECT 101.530 10.090 101.790 11.225 ;
        RECT 101.980 10.295 102.210 11.605 ;
        RECT 102.755 11.545 103.015 11.865 ;
        RECT 103.345 11.545 103.605 11.865 ;
        RECT 104.135 11.545 104.395 11.865 ;
        RECT 102.770 10.295 103.000 11.545 ;
        RECT 103.360 10.295 103.590 11.545 ;
        RECT 104.150 10.295 104.380 11.545 ;
        RECT 104.620 10.090 104.880 10.595 ;
        RECT 101.530 9.860 102.720 10.090 ;
        RECT 103.640 9.860 104.880 10.090 ;
        RECT 105.305 10.230 105.660 11.835 ;
        RECT 106.040 10.230 106.395 11.840 ;
        RECT 107.315 11.775 107.545 12.740 ;
        RECT 108.105 11.865 108.335 12.740 ;
        RECT 108.695 11.865 108.925 12.740 ;
        RECT 109.485 11.865 109.715 12.740 ;
        RECT 109.955 12.110 110.215 12.900 ;
        RECT 112.140 12.900 113.380 13.130 ;
        RECT 114.300 12.900 115.540 13.130 ;
        RECT 112.140 12.205 112.400 12.900 ;
        RECT 105.305 9.645 106.395 10.230 ;
        RECT 106.535 11.605 107.545 11.775 ;
        RECT 106.535 9.645 106.705 11.605 ;
        RECT 106.865 10.090 107.125 11.225 ;
        RECT 107.315 10.295 107.545 11.605 ;
        RECT 108.090 11.545 108.350 11.865 ;
        RECT 108.680 11.545 108.940 11.865 ;
        RECT 109.470 11.545 109.730 11.865 ;
        RECT 108.105 10.295 108.335 11.545 ;
        RECT 108.695 10.295 108.925 11.545 ;
        RECT 109.485 10.295 109.715 11.545 ;
        RECT 109.955 10.090 110.215 10.595 ;
        RECT 106.865 9.860 108.055 10.090 ;
        RECT 108.975 9.860 110.215 10.090 ;
        RECT 110.640 10.235 110.995 11.835 ;
        RECT 111.365 10.235 111.720 11.840 ;
        RECT 112.640 11.775 112.870 12.740 ;
        RECT 113.430 11.865 113.660 12.740 ;
        RECT 114.020 11.865 114.250 12.740 ;
        RECT 114.810 11.865 115.040 12.740 ;
        RECT 115.280 12.110 115.540 12.900 ;
        RECT 117.475 12.900 118.715 13.130 ;
        RECT 119.635 12.900 120.875 13.130 ;
        RECT 117.475 12.205 117.735 12.900 ;
        RECT 110.640 9.650 111.720 10.235 ;
        RECT 110.640 9.645 110.995 9.650 ;
        RECT 100.705 9.370 101.370 9.645 ;
        RECT 104.990 9.370 105.660 9.645 ;
        RECT 100.705 7.265 101.060 9.370 ;
        RECT 101.980 7.505 102.210 8.740 ;
        RECT 102.770 7.505 103.000 8.740 ;
        RECT 103.360 7.505 103.590 8.740 ;
        RECT 96.655 6.295 96.885 7.185 ;
        RECT 97.445 6.295 97.675 7.185 ;
        RECT 98.035 6.295 98.265 7.185 ;
        RECT 98.825 6.295 99.055 7.260 ;
        RECT 101.965 7.185 102.225 7.505 ;
        RECT 102.755 7.185 103.015 7.505 ;
        RECT 103.345 7.185 103.605 7.505 ;
        RECT 104.150 7.430 104.380 8.740 ;
        RECT 104.990 7.430 105.160 9.370 ;
        RECT 104.150 7.260 105.160 7.430 ;
        RECT 105.305 7.260 105.660 9.370 ;
        RECT 106.040 9.370 106.705 9.645 ;
        RECT 110.325 9.370 110.995 9.645 ;
        RECT 106.040 7.265 106.395 9.370 ;
        RECT 107.315 7.505 107.545 8.740 ;
        RECT 108.105 7.505 108.335 8.740 ;
        RECT 108.695 7.505 108.925 8.740 ;
        RECT 101.980 6.295 102.210 7.185 ;
        RECT 102.770 6.295 103.000 7.185 ;
        RECT 103.360 6.295 103.590 7.185 ;
        RECT 104.150 6.295 104.380 7.260 ;
        RECT 107.300 7.185 107.560 7.505 ;
        RECT 108.090 7.185 108.350 7.505 ;
        RECT 108.680 7.185 108.940 7.505 ;
        RECT 109.485 7.430 109.715 8.740 ;
        RECT 110.325 7.430 110.495 9.370 ;
        RECT 109.485 7.260 110.495 7.430 ;
        RECT 110.640 7.260 110.995 9.370 ;
        RECT 111.365 9.645 111.720 9.650 ;
        RECT 111.860 11.605 112.870 11.775 ;
        RECT 111.860 9.645 112.030 11.605 ;
        RECT 112.190 10.090 112.450 11.225 ;
        RECT 112.640 10.295 112.870 11.605 ;
        RECT 113.415 11.545 113.675 11.865 ;
        RECT 114.005 11.545 114.265 11.865 ;
        RECT 114.795 11.545 115.055 11.865 ;
        RECT 113.430 10.295 113.660 11.545 ;
        RECT 114.020 10.295 114.250 11.545 ;
        RECT 114.810 10.295 115.040 11.545 ;
        RECT 115.280 10.090 115.540 10.595 ;
        RECT 112.190 9.860 113.380 10.090 ;
        RECT 114.300 9.860 115.540 10.090 ;
        RECT 115.965 10.230 116.320 11.835 ;
        RECT 116.700 10.230 117.055 11.840 ;
        RECT 117.975 11.775 118.205 12.740 ;
        RECT 118.765 11.865 118.995 12.740 ;
        RECT 119.355 11.865 119.585 12.740 ;
        RECT 120.145 11.865 120.375 12.740 ;
        RECT 120.615 12.110 120.875 12.900 ;
        RECT 124.090 11.865 124.320 12.740 ;
        RECT 124.680 11.865 124.910 12.740 ;
        RECT 125.470 11.865 125.700 12.740 ;
        RECT 115.965 9.645 117.055 10.230 ;
        RECT 117.195 11.605 118.205 11.775 ;
        RECT 117.195 9.645 117.365 11.605 ;
        RECT 117.525 10.090 117.785 11.225 ;
        RECT 117.975 10.295 118.205 11.605 ;
        RECT 118.750 11.545 119.010 11.865 ;
        RECT 119.340 11.545 119.600 11.865 ;
        RECT 120.130 11.545 120.390 11.865 ;
        RECT 124.075 11.545 124.335 11.865 ;
        RECT 124.665 11.545 124.925 11.865 ;
        RECT 125.455 11.545 125.715 11.865 ;
        RECT 118.765 10.295 118.995 11.545 ;
        RECT 119.355 10.295 119.585 11.545 ;
        RECT 120.145 10.295 120.375 11.545 ;
        RECT 120.615 10.090 120.875 10.595 ;
        RECT 124.090 10.295 124.320 11.545 ;
        RECT 124.680 10.295 124.910 11.545 ;
        RECT 125.470 10.295 125.700 11.545 ;
        RECT 117.525 9.860 118.715 10.090 ;
        RECT 119.635 9.860 120.875 10.090 ;
        RECT 126.625 10.235 126.980 11.855 ;
        RECT 126.625 9.650 127.170 10.235 ;
        RECT 126.625 9.645 126.980 9.650 ;
        RECT 111.365 9.370 112.030 9.645 ;
        RECT 115.650 9.370 116.320 9.645 ;
        RECT 111.365 7.265 111.720 9.370 ;
        RECT 112.640 7.505 112.870 8.740 ;
        RECT 113.430 7.505 113.660 8.740 ;
        RECT 114.020 7.505 114.250 8.740 ;
        RECT 107.315 6.295 107.545 7.185 ;
        RECT 108.105 6.295 108.335 7.185 ;
        RECT 108.695 6.295 108.925 7.185 ;
        RECT 109.485 6.295 109.715 7.260 ;
        RECT 112.625 7.185 112.885 7.505 ;
        RECT 113.415 7.185 113.675 7.505 ;
        RECT 114.005 7.185 114.265 7.505 ;
        RECT 114.810 7.430 115.040 8.740 ;
        RECT 115.650 7.430 115.820 9.370 ;
        RECT 114.810 7.260 115.820 7.430 ;
        RECT 115.965 7.260 116.320 9.370 ;
        RECT 116.700 9.370 117.365 9.645 ;
        RECT 126.310 9.370 126.980 9.645 ;
        RECT 116.700 7.265 117.055 9.370 ;
        RECT 117.975 7.505 118.205 8.740 ;
        RECT 118.765 7.505 118.995 8.740 ;
        RECT 119.355 7.505 119.585 8.740 ;
        RECT 123.300 7.505 123.530 8.740 ;
        RECT 124.090 7.505 124.320 8.740 ;
        RECT 124.680 7.505 124.910 8.740 ;
        RECT 112.640 6.295 112.870 7.185 ;
        RECT 113.430 6.295 113.660 7.185 ;
        RECT 114.020 6.295 114.250 7.185 ;
        RECT 114.810 6.295 115.040 7.260 ;
        RECT 117.960 7.185 118.220 7.505 ;
        RECT 118.750 7.185 119.010 7.505 ;
        RECT 119.340 7.185 119.600 7.505 ;
        RECT 123.285 7.185 123.545 7.505 ;
        RECT 124.075 7.185 124.335 7.505 ;
        RECT 124.665 7.185 124.925 7.505 ;
        RECT 125.470 7.430 125.700 8.740 ;
        RECT 126.310 7.430 126.480 9.370 ;
        RECT 125.470 7.260 126.480 7.430 ;
        RECT 126.625 7.280 126.980 9.370 ;
        RECT 117.975 6.295 118.205 7.185 ;
        RECT 118.765 6.295 118.995 7.185 ;
        RECT 119.355 6.295 119.585 7.185 ;
        RECT 123.300 6.295 123.530 7.185 ;
        RECT 124.090 6.295 124.320 7.185 ;
        RECT 124.680 6.295 124.910 7.185 ;
        RECT 125.470 6.295 125.700 7.260 ;
        RECT 10.500 3.630 10.820 4.115 ;
        RECT 16.115 3.740 28.735 3.975 ;
        RECT 10.500 3.300 11.960 3.630 ;
        RECT 10.500 3.080 10.820 3.300 ;
        RECT 12.400 2.555 12.720 3.545 ;
        RECT 14.585 3.300 16.005 3.625 ;
        RECT 19.990 3.170 28.735 3.740 ;
        RECT 16.115 2.935 28.735 3.170 ;
        RECT 12.425 2.540 12.715 2.555 ;
        RECT 31.420 2.110 31.775 4.320 ;
        RECT 32.695 4.240 32.925 5.205 ;
        RECT 33.485 4.330 33.715 5.205 ;
        RECT 34.075 4.330 34.305 5.205 ;
        RECT 34.865 4.330 35.095 5.205 ;
        RECT 31.915 4.070 32.925 4.240 ;
        RECT 31.915 2.110 32.085 4.070 ;
        RECT 32.695 2.760 32.925 4.070 ;
        RECT 33.470 4.010 33.730 4.330 ;
        RECT 34.060 4.010 34.320 4.330 ;
        RECT 34.850 4.010 35.110 4.330 ;
        RECT 33.485 2.760 33.715 4.010 ;
        RECT 34.075 2.760 34.305 4.010 ;
        RECT 34.865 2.760 35.095 4.010 ;
        RECT 31.240 1.835 32.085 2.110 ;
        RECT 36.020 2.110 36.375 4.320 ;
        RECT 36.745 2.110 37.100 4.305 ;
        RECT 38.020 4.240 38.250 5.205 ;
        RECT 38.810 4.330 39.040 5.205 ;
        RECT 39.400 4.330 39.630 5.205 ;
        RECT 40.190 4.330 40.420 5.205 ;
        RECT 37.240 4.070 38.250 4.240 ;
        RECT 37.240 2.110 37.410 4.070 ;
        RECT 38.020 2.760 38.250 4.070 ;
        RECT 38.795 4.010 39.055 4.330 ;
        RECT 39.385 4.010 39.645 4.330 ;
        RECT 40.175 4.010 40.435 4.330 ;
        RECT 38.810 2.760 39.040 4.010 ;
        RECT 39.400 2.760 39.630 4.010 ;
        RECT 40.190 2.760 40.420 4.010 ;
        RECT 36.020 1.835 37.410 2.110 ;
        RECT 41.345 2.110 41.700 4.300 ;
        RECT 42.080 2.110 42.435 4.305 ;
        RECT 43.355 4.240 43.585 5.205 ;
        RECT 44.145 4.330 44.375 5.205 ;
        RECT 44.735 4.330 44.965 5.205 ;
        RECT 45.525 4.330 45.755 5.205 ;
        RECT 42.575 4.070 43.585 4.240 ;
        RECT 42.575 2.110 42.745 4.070 ;
        RECT 43.355 2.760 43.585 4.070 ;
        RECT 44.130 4.010 44.390 4.330 ;
        RECT 44.720 4.010 44.980 4.330 ;
        RECT 45.510 4.010 45.770 4.330 ;
        RECT 44.145 2.760 44.375 4.010 ;
        RECT 44.735 2.760 44.965 4.010 ;
        RECT 45.525 2.760 45.755 4.010 ;
        RECT 41.345 1.835 42.745 2.110 ;
        RECT 46.680 2.110 47.035 4.300 ;
        RECT 47.405 2.110 47.760 4.305 ;
        RECT 48.680 4.240 48.910 5.205 ;
        RECT 49.470 4.330 49.700 5.205 ;
        RECT 50.060 4.330 50.290 5.205 ;
        RECT 50.850 4.330 51.080 5.205 ;
        RECT 47.900 4.070 48.910 4.240 ;
        RECT 47.900 2.110 48.070 4.070 ;
        RECT 48.680 2.760 48.910 4.070 ;
        RECT 49.455 4.010 49.715 4.330 ;
        RECT 50.045 4.010 50.305 4.330 ;
        RECT 50.835 4.010 51.095 4.330 ;
        RECT 49.470 2.760 49.700 4.010 ;
        RECT 50.060 2.760 50.290 4.010 ;
        RECT 50.850 2.760 51.080 4.010 ;
        RECT 46.680 1.835 48.070 2.110 ;
        RECT 52.005 2.110 52.360 4.300 ;
        RECT 52.740 2.110 53.095 4.305 ;
        RECT 54.015 4.240 54.245 5.205 ;
        RECT 54.805 4.330 55.035 5.205 ;
        RECT 55.395 4.330 55.625 5.205 ;
        RECT 56.185 4.330 56.415 5.205 ;
        RECT 53.235 4.070 54.245 4.240 ;
        RECT 53.235 2.110 53.405 4.070 ;
        RECT 54.015 2.760 54.245 4.070 ;
        RECT 54.790 4.010 55.050 4.330 ;
        RECT 55.380 4.010 55.640 4.330 ;
        RECT 56.170 4.010 56.430 4.330 ;
        RECT 54.805 2.760 55.035 4.010 ;
        RECT 55.395 2.760 55.625 4.010 ;
        RECT 56.185 2.760 56.415 4.010 ;
        RECT 52.005 1.835 53.405 2.110 ;
        RECT 57.340 2.110 57.695 4.300 ;
        RECT 58.065 2.110 58.420 4.305 ;
        RECT 59.340 4.240 59.570 5.205 ;
        RECT 60.130 4.330 60.360 5.205 ;
        RECT 60.720 4.330 60.950 5.205 ;
        RECT 61.510 4.330 61.740 5.205 ;
        RECT 58.560 4.070 59.570 4.240 ;
        RECT 58.560 2.110 58.730 4.070 ;
        RECT 59.340 2.760 59.570 4.070 ;
        RECT 60.115 4.010 60.375 4.330 ;
        RECT 60.705 4.010 60.965 4.330 ;
        RECT 61.495 4.010 61.755 4.330 ;
        RECT 60.130 2.760 60.360 4.010 ;
        RECT 60.720 2.760 60.950 4.010 ;
        RECT 61.510 2.760 61.740 4.010 ;
        RECT 57.340 1.835 58.730 2.110 ;
        RECT 62.665 2.110 63.020 4.300 ;
        RECT 63.400 2.110 63.755 4.305 ;
        RECT 64.675 4.240 64.905 5.205 ;
        RECT 65.465 4.330 65.695 5.205 ;
        RECT 66.055 4.330 66.285 5.205 ;
        RECT 66.845 4.330 67.075 5.205 ;
        RECT 63.895 4.070 64.905 4.240 ;
        RECT 63.895 2.110 64.065 4.070 ;
        RECT 64.675 2.760 64.905 4.070 ;
        RECT 65.450 4.010 65.710 4.330 ;
        RECT 66.040 4.010 66.300 4.330 ;
        RECT 66.830 4.010 67.090 4.330 ;
        RECT 65.465 2.760 65.695 4.010 ;
        RECT 66.055 2.760 66.285 4.010 ;
        RECT 66.845 2.760 67.075 4.010 ;
        RECT 62.665 1.835 64.065 2.110 ;
        RECT 68.000 2.110 68.355 4.300 ;
        RECT 68.725 2.110 69.080 4.305 ;
        RECT 70.000 4.240 70.230 5.205 ;
        RECT 70.790 4.330 71.020 5.205 ;
        RECT 71.380 4.330 71.610 5.205 ;
        RECT 72.170 4.330 72.400 5.205 ;
        RECT 69.220 4.070 70.230 4.240 ;
        RECT 69.220 2.110 69.390 4.070 ;
        RECT 70.000 2.760 70.230 4.070 ;
        RECT 70.775 4.010 71.035 4.330 ;
        RECT 71.365 4.010 71.625 4.330 ;
        RECT 72.155 4.010 72.415 4.330 ;
        RECT 70.790 2.760 71.020 4.010 ;
        RECT 71.380 2.760 71.610 4.010 ;
        RECT 72.170 2.760 72.400 4.010 ;
        RECT 68.000 1.835 69.390 2.110 ;
        RECT 73.325 2.110 73.680 4.300 ;
        RECT 74.060 2.110 74.415 4.305 ;
        RECT 75.335 4.240 75.565 5.205 ;
        RECT 76.125 4.330 76.355 5.205 ;
        RECT 76.715 4.330 76.945 5.205 ;
        RECT 77.505 4.330 77.735 5.205 ;
        RECT 74.555 4.070 75.565 4.240 ;
        RECT 74.555 2.110 74.725 4.070 ;
        RECT 75.335 2.760 75.565 4.070 ;
        RECT 76.110 4.010 76.370 4.330 ;
        RECT 76.700 4.010 76.960 4.330 ;
        RECT 77.490 4.010 77.750 4.330 ;
        RECT 76.125 2.760 76.355 4.010 ;
        RECT 76.715 2.760 76.945 4.010 ;
        RECT 77.505 2.760 77.735 4.010 ;
        RECT 73.325 1.835 74.725 2.110 ;
        RECT 78.660 2.110 79.015 4.300 ;
        RECT 79.385 2.110 79.740 4.305 ;
        RECT 80.660 4.240 80.890 5.205 ;
        RECT 81.450 4.330 81.680 5.205 ;
        RECT 82.040 4.330 82.270 5.205 ;
        RECT 82.830 4.330 83.060 5.205 ;
        RECT 79.880 4.070 80.890 4.240 ;
        RECT 79.880 2.110 80.050 4.070 ;
        RECT 80.660 2.760 80.890 4.070 ;
        RECT 81.435 4.010 81.695 4.330 ;
        RECT 82.025 4.010 82.285 4.330 ;
        RECT 82.815 4.010 83.075 4.330 ;
        RECT 81.450 2.760 81.680 4.010 ;
        RECT 82.040 2.760 82.270 4.010 ;
        RECT 82.830 2.760 83.060 4.010 ;
        RECT 78.660 1.835 80.050 2.110 ;
        RECT 83.985 2.110 84.340 4.300 ;
        RECT 84.720 2.110 85.075 4.305 ;
        RECT 85.995 4.240 86.225 5.205 ;
        RECT 86.785 4.330 87.015 5.205 ;
        RECT 87.375 4.330 87.605 5.205 ;
        RECT 88.165 4.330 88.395 5.205 ;
        RECT 85.215 4.070 86.225 4.240 ;
        RECT 85.215 2.110 85.385 4.070 ;
        RECT 85.995 2.760 86.225 4.070 ;
        RECT 86.770 4.010 87.030 4.330 ;
        RECT 87.360 4.010 87.620 4.330 ;
        RECT 88.150 4.010 88.410 4.330 ;
        RECT 86.785 2.760 87.015 4.010 ;
        RECT 87.375 2.760 87.605 4.010 ;
        RECT 88.165 2.760 88.395 4.010 ;
        RECT 83.985 1.835 85.385 2.110 ;
        RECT 89.320 2.110 89.675 4.300 ;
        RECT 90.045 2.110 90.400 4.305 ;
        RECT 91.320 4.240 91.550 5.205 ;
        RECT 92.110 4.330 92.340 5.205 ;
        RECT 92.700 4.330 92.930 5.205 ;
        RECT 93.490 4.330 93.720 5.205 ;
        RECT 90.540 4.070 91.550 4.240 ;
        RECT 90.540 2.110 90.710 4.070 ;
        RECT 91.320 2.760 91.550 4.070 ;
        RECT 92.095 4.010 92.355 4.330 ;
        RECT 92.685 4.010 92.945 4.330 ;
        RECT 93.475 4.010 93.735 4.330 ;
        RECT 92.110 2.760 92.340 4.010 ;
        RECT 92.700 2.760 92.930 4.010 ;
        RECT 93.490 2.760 93.720 4.010 ;
        RECT 89.320 1.835 90.710 2.110 ;
        RECT 94.645 2.110 95.000 4.300 ;
        RECT 95.380 2.110 95.735 4.305 ;
        RECT 96.655 4.240 96.885 5.205 ;
        RECT 97.445 4.330 97.675 5.205 ;
        RECT 98.035 4.330 98.265 5.205 ;
        RECT 98.825 4.330 99.055 5.205 ;
        RECT 95.875 4.070 96.885 4.240 ;
        RECT 95.875 2.110 96.045 4.070 ;
        RECT 96.655 2.760 96.885 4.070 ;
        RECT 97.430 4.010 97.690 4.330 ;
        RECT 98.020 4.010 98.280 4.330 ;
        RECT 98.810 4.010 99.070 4.330 ;
        RECT 97.445 2.760 97.675 4.010 ;
        RECT 98.035 2.760 98.265 4.010 ;
        RECT 98.825 2.760 99.055 4.010 ;
        RECT 94.645 1.835 96.045 2.110 ;
        RECT 99.980 2.110 100.335 4.300 ;
        RECT 100.705 2.110 101.060 4.305 ;
        RECT 101.980 4.240 102.210 5.205 ;
        RECT 102.770 4.330 103.000 5.205 ;
        RECT 103.360 4.330 103.590 5.205 ;
        RECT 104.150 4.330 104.380 5.205 ;
        RECT 101.200 4.070 102.210 4.240 ;
        RECT 101.200 2.110 101.370 4.070 ;
        RECT 101.980 2.760 102.210 4.070 ;
        RECT 102.755 4.010 103.015 4.330 ;
        RECT 103.345 4.010 103.605 4.330 ;
        RECT 104.135 4.010 104.395 4.330 ;
        RECT 102.770 2.760 103.000 4.010 ;
        RECT 103.360 2.760 103.590 4.010 ;
        RECT 104.150 2.760 104.380 4.010 ;
        RECT 99.980 1.835 101.370 2.110 ;
        RECT 105.305 2.110 105.660 4.300 ;
        RECT 106.040 2.110 106.395 4.305 ;
        RECT 107.315 4.240 107.545 5.205 ;
        RECT 108.105 4.330 108.335 5.205 ;
        RECT 108.695 4.330 108.925 5.205 ;
        RECT 109.485 4.330 109.715 5.205 ;
        RECT 106.535 4.070 107.545 4.240 ;
        RECT 106.535 2.110 106.705 4.070 ;
        RECT 107.315 2.760 107.545 4.070 ;
        RECT 108.090 4.010 108.350 4.330 ;
        RECT 108.680 4.010 108.940 4.330 ;
        RECT 109.470 4.010 109.730 4.330 ;
        RECT 108.105 2.760 108.335 4.010 ;
        RECT 108.695 2.760 108.925 4.010 ;
        RECT 109.485 2.760 109.715 4.010 ;
        RECT 105.305 1.835 106.705 2.110 ;
        RECT 110.640 2.110 110.995 4.300 ;
        RECT 111.365 2.110 111.720 4.305 ;
        RECT 112.640 4.240 112.870 5.205 ;
        RECT 113.430 4.330 113.660 5.205 ;
        RECT 114.020 4.330 114.250 5.205 ;
        RECT 114.810 4.330 115.040 5.205 ;
        RECT 111.860 4.070 112.870 4.240 ;
        RECT 111.860 2.110 112.030 4.070 ;
        RECT 112.640 2.760 112.870 4.070 ;
        RECT 113.415 4.010 113.675 4.330 ;
        RECT 114.005 4.010 114.265 4.330 ;
        RECT 114.795 4.010 115.055 4.330 ;
        RECT 113.430 2.760 113.660 4.010 ;
        RECT 114.020 2.760 114.250 4.010 ;
        RECT 114.810 2.760 115.040 4.010 ;
        RECT 110.640 1.835 112.030 2.110 ;
        RECT 115.965 2.110 116.320 4.300 ;
        RECT 116.700 2.110 117.055 4.305 ;
        RECT 117.975 4.240 118.205 5.205 ;
        RECT 118.765 4.330 118.995 5.205 ;
        RECT 119.355 4.330 119.585 5.205 ;
        RECT 120.145 4.330 120.375 5.205 ;
        RECT 117.195 4.070 118.205 4.240 ;
        RECT 117.195 2.110 117.365 4.070 ;
        RECT 117.975 2.760 118.205 4.070 ;
        RECT 118.750 4.010 119.010 4.330 ;
        RECT 119.340 4.010 119.600 4.330 ;
        RECT 120.130 4.010 120.390 4.330 ;
        RECT 118.765 2.760 118.995 4.010 ;
        RECT 119.355 2.760 119.585 4.010 ;
        RECT 120.145 2.760 120.375 4.010 ;
        RECT 115.965 1.835 117.365 2.110 ;
        RECT 121.300 2.110 121.655 4.300 ;
        RECT 122.025 2.110 122.380 4.320 ;
        RECT 123.300 4.240 123.530 5.205 ;
        RECT 124.090 4.330 124.320 5.205 ;
        RECT 124.680 4.330 124.910 5.205 ;
        RECT 125.470 4.330 125.700 5.205 ;
        RECT 122.520 4.070 123.530 4.240 ;
        RECT 122.520 2.110 122.690 4.070 ;
        RECT 123.300 2.760 123.530 4.070 ;
        RECT 124.075 4.010 124.335 4.330 ;
        RECT 124.665 4.010 124.925 4.330 ;
        RECT 125.455 4.010 125.715 4.330 ;
        RECT 126.685 4.320 126.935 7.280 ;
        RECT 124.090 2.760 124.320 4.010 ;
        RECT 124.680 2.760 124.910 4.010 ;
        RECT 125.470 2.760 125.700 4.010 ;
        RECT 121.300 1.835 122.690 2.110 ;
        RECT 126.625 2.110 126.980 4.320 ;
        RECT 126.625 1.835 127.170 2.110 ;
      LAYER met2 ;
        RECT 53.435 80.775 53.805 80.825 ;
        RECT 96.705 80.775 97.075 80.830 ;
        RECT 22.765 80.595 97.085 80.775 ;
        RECT 22.765 65.715 22.945 80.595 ;
        RECT 53.435 80.545 53.805 80.595 ;
        RECT 96.705 80.550 97.075 80.595 ;
        RECT 54.065 80.395 54.435 80.435 ;
        RECT 96.075 80.395 96.445 80.445 ;
        RECT 23.145 80.215 96.485 80.395 ;
        RECT 10.530 60.060 10.790 65.575 ;
        RECT 11.745 65.055 13.345 65.345 ;
        RECT 12.430 59.505 12.690 65.055 ;
        RECT 16.040 64.610 17.645 64.900 ;
        RECT 16.110 64.050 16.565 64.610 ;
        RECT 22.725 64.605 22.985 65.715 ;
        RECT 22.765 64.580 22.945 64.605 ;
        RECT 15.455 63.595 16.565 64.050 ;
        RECT 15.455 60.590 15.910 63.595 ;
        RECT 23.145 60.985 23.325 80.215 ;
        RECT 54.065 80.155 54.435 80.215 ;
        RECT 96.075 80.165 96.445 80.215 ;
        RECT 42.775 80.015 43.145 80.065 ;
        RECT 64.725 80.015 65.095 80.055 ;
        RECT 85.415 80.015 85.785 80.065 ;
        RECT 107.365 80.015 107.735 80.055 ;
        RECT 23.525 79.835 107.760 80.015 ;
        RECT 14.605 60.300 15.985 60.590 ;
        RECT 23.105 59.880 23.365 60.985 ;
        RECT 23.145 59.805 23.325 59.880 ;
        RECT 23.525 57.575 23.705 79.835 ;
        RECT 42.775 79.785 43.145 79.835 ;
        RECT 64.725 79.775 65.095 79.835 ;
        RECT 85.415 79.785 85.785 79.835 ;
        RECT 107.365 79.775 107.735 79.835 ;
        RECT 43.405 79.635 43.775 79.675 ;
        RECT 64.095 79.635 64.465 79.685 ;
        RECT 86.045 79.635 86.415 79.675 ;
        RECT 106.735 79.635 107.105 79.685 ;
        RECT 23.905 79.455 107.155 79.635 ;
        RECT 10.530 51.920 10.790 57.435 ;
        RECT 11.745 56.915 13.345 57.205 ;
        RECT 12.430 51.365 12.690 56.915 ;
        RECT 16.040 56.470 17.645 56.760 ;
        RECT 16.110 55.910 16.565 56.470 ;
        RECT 23.485 56.465 23.745 57.575 ;
        RECT 23.525 56.410 23.705 56.465 ;
        RECT 15.455 55.455 16.565 55.910 ;
        RECT 15.455 52.450 15.910 55.455 ;
        RECT 23.905 52.850 24.085 79.455 ;
        RECT 43.405 79.395 43.775 79.455 ;
        RECT 64.095 79.405 64.465 79.455 ;
        RECT 86.045 79.395 86.415 79.455 ;
        RECT 106.735 79.405 107.105 79.455 ;
        RECT 32.625 75.020 34.390 75.300 ;
        RECT 37.950 75.020 39.715 75.300 ;
        RECT 43.285 75.020 45.050 75.300 ;
        RECT 48.610 75.020 50.375 75.300 ;
        RECT 53.945 75.020 55.710 75.300 ;
        RECT 59.270 75.020 61.035 75.300 ;
        RECT 64.605 75.020 66.370 75.300 ;
        RECT 69.930 75.020 71.695 75.300 ;
        RECT 75.265 75.020 77.030 75.300 ;
        RECT 80.590 75.020 82.355 75.300 ;
        RECT 85.925 75.020 87.690 75.300 ;
        RECT 91.250 75.020 93.015 75.300 ;
        RECT 96.585 75.020 98.350 75.300 ;
        RECT 101.910 75.020 103.675 75.300 ;
        RECT 107.245 75.020 109.010 75.300 ;
        RECT 112.570 75.020 114.335 75.300 ;
        RECT 117.905 75.020 119.670 75.300 ;
        RECT 123.230 75.020 124.995 75.300 ;
        RECT 34.005 72.125 34.400 72.130 ;
        RECT 38.900 72.125 40.145 72.130 ;
        RECT 44.280 72.125 45.470 72.130 ;
        RECT 49.560 72.125 50.805 72.130 ;
        RECT 54.940 72.125 56.130 72.130 ;
        RECT 60.220 72.125 61.465 72.130 ;
        RECT 65.600 72.125 66.790 72.130 ;
        RECT 70.880 72.125 72.125 72.130 ;
        RECT 76.260 72.125 77.450 72.130 ;
        RECT 81.540 72.125 82.785 72.130 ;
        RECT 86.920 72.125 88.110 72.130 ;
        RECT 92.200 72.125 93.445 72.130 ;
        RECT 97.580 72.125 98.770 72.130 ;
        RECT 102.860 72.125 104.105 72.130 ;
        RECT 108.240 72.125 109.430 72.130 ;
        RECT 113.520 72.125 114.765 72.130 ;
        RECT 118.900 72.125 120.090 72.130 ;
        RECT 124.610 72.125 125.005 72.130 ;
        RECT 33.390 71.845 35.160 72.125 ;
        RECT 38.715 71.850 40.485 72.125 ;
        RECT 38.715 71.845 39.110 71.850 ;
        RECT 40.120 71.845 40.485 71.850 ;
        RECT 44.050 71.850 45.820 72.125 ;
        RECT 44.050 71.845 44.445 71.850 ;
        RECT 45.455 71.845 45.820 71.850 ;
        RECT 49.375 71.850 51.145 72.125 ;
        RECT 49.375 71.845 49.770 71.850 ;
        RECT 50.780 71.845 51.145 71.850 ;
        RECT 54.710 71.850 56.480 72.125 ;
        RECT 54.710 71.845 55.105 71.850 ;
        RECT 56.115 71.845 56.480 71.850 ;
        RECT 60.035 71.850 61.805 72.125 ;
        RECT 60.035 71.845 60.430 71.850 ;
        RECT 61.440 71.845 61.805 71.850 ;
        RECT 65.370 71.850 67.140 72.125 ;
        RECT 65.370 71.845 65.765 71.850 ;
        RECT 66.775 71.845 67.140 71.850 ;
        RECT 70.695 71.850 72.465 72.125 ;
        RECT 70.695 71.845 71.090 71.850 ;
        RECT 72.100 71.845 72.465 71.850 ;
        RECT 76.030 71.850 77.800 72.125 ;
        RECT 76.030 71.845 76.425 71.850 ;
        RECT 77.435 71.845 77.800 71.850 ;
        RECT 81.355 71.850 83.125 72.125 ;
        RECT 81.355 71.845 81.750 71.850 ;
        RECT 82.760 71.845 83.125 71.850 ;
        RECT 86.690 71.850 88.460 72.125 ;
        RECT 86.690 71.845 87.085 71.850 ;
        RECT 88.095 71.845 88.460 71.850 ;
        RECT 92.015 71.850 93.785 72.125 ;
        RECT 92.015 71.845 92.410 71.850 ;
        RECT 93.420 71.845 93.785 71.850 ;
        RECT 97.350 71.850 99.120 72.125 ;
        RECT 97.350 71.845 97.745 71.850 ;
        RECT 98.755 71.845 99.120 71.850 ;
        RECT 102.675 71.850 104.445 72.125 ;
        RECT 102.675 71.845 103.070 71.850 ;
        RECT 104.080 71.845 104.445 71.850 ;
        RECT 108.010 71.850 109.780 72.125 ;
        RECT 108.010 71.845 108.405 71.850 ;
        RECT 109.415 71.845 109.780 71.850 ;
        RECT 113.335 71.850 115.105 72.125 ;
        RECT 113.335 71.845 113.730 71.850 ;
        RECT 114.740 71.845 115.105 71.850 ;
        RECT 118.670 71.850 120.440 72.125 ;
        RECT 118.670 71.845 119.065 71.850 ;
        RECT 120.075 71.845 120.440 71.850 ;
        RECT 123.995 71.845 125.765 72.125 ;
        RECT 24.285 67.570 24.465 69.890 ;
        RECT 24.665 68.860 24.845 69.890 ;
        RECT 24.610 68.490 24.890 68.860 ;
        RECT 24.235 67.200 24.515 67.570 ;
        RECT 14.605 52.160 15.985 52.450 ;
        RECT 23.865 51.745 24.125 52.850 ;
        RECT 23.905 51.700 24.085 51.745 ;
        RECT 10.530 43.780 10.790 49.295 ;
        RECT 11.745 48.775 13.345 49.065 ;
        RECT 12.430 43.225 12.690 48.775 ;
        RECT 16.040 48.330 17.645 48.620 ;
        RECT 16.110 47.770 16.565 48.330 ;
        RECT 15.455 47.315 16.565 47.770 ;
        RECT 15.455 44.310 15.910 47.315 ;
        RECT 24.285 44.710 24.465 67.200 ;
        RECT 24.665 49.435 24.845 68.490 ;
        RECT 24.625 48.325 24.885 49.435 ;
        RECT 24.665 48.310 24.845 48.325 ;
        RECT 14.605 44.020 15.985 44.310 ;
        RECT 24.245 43.605 24.505 44.710 ;
        RECT 24.285 43.550 24.465 43.605 ;
        RECT 10.530 35.640 10.790 41.155 ;
        RECT 11.745 40.635 13.345 40.925 ;
        RECT 12.430 35.085 12.690 40.635 ;
        RECT 16.040 40.190 17.645 40.480 ;
        RECT 16.110 39.630 16.565 40.190 ;
        RECT 15.455 39.175 16.565 39.630 ;
        RECT 15.455 36.170 15.910 39.175 ;
        RECT 25.045 36.570 25.225 69.890 ;
        RECT 25.425 40.295 25.605 69.890 ;
        RECT 25.805 41.050 25.985 69.890 ;
        RECT 26.185 42.340 26.365 69.890 ;
        RECT 26.565 57.410 26.745 69.890 ;
        RECT 26.515 57.040 26.795 57.410 ;
        RECT 26.565 53.790 26.745 57.040 ;
        RECT 26.945 56.120 27.125 69.890 ;
        RECT 27.325 64.945 27.505 69.890 ;
        RECT 27.275 64.575 27.555 64.945 ;
        RECT 27.325 61.325 27.505 64.575 ;
        RECT 27.705 63.655 27.885 69.890 ;
        RECT 28.085 68.215 28.265 69.890 ;
        RECT 28.035 67.845 28.315 68.215 ;
        RECT 28.085 65.595 28.265 67.845 ;
        RECT 28.465 66.925 28.645 69.890 ;
        RECT 36.790 69.110 37.160 69.120 ;
        RECT 36.790 68.850 37.810 69.110 ;
        RECT 40.960 68.930 41.600 69.140 ;
        RECT 36.790 68.840 37.160 68.850 ;
        RECT 39.895 68.810 41.600 68.930 ;
        RECT 42.125 69.110 42.495 69.120 ;
        RECT 42.125 68.850 43.145 69.110 ;
        RECT 46.295 68.930 46.935 69.140 ;
        RECT 42.125 68.840 42.495 68.850 ;
        RECT 45.230 68.810 46.935 68.930 ;
        RECT 47.450 69.110 47.820 69.120 ;
        RECT 47.450 68.850 48.470 69.110 ;
        RECT 51.620 68.930 52.260 69.140 ;
        RECT 47.450 68.840 47.820 68.850 ;
        RECT 50.555 68.810 52.260 68.930 ;
        RECT 52.785 69.110 53.155 69.120 ;
        RECT 52.785 68.850 53.805 69.110 ;
        RECT 56.955 68.930 57.595 69.140 ;
        RECT 52.785 68.840 53.155 68.850 ;
        RECT 55.890 68.810 57.595 68.930 ;
        RECT 58.110 69.110 58.480 69.120 ;
        RECT 58.110 68.850 59.130 69.110 ;
        RECT 62.280 68.930 62.920 69.140 ;
        RECT 58.110 68.840 58.480 68.850 ;
        RECT 61.215 68.810 62.920 68.930 ;
        RECT 63.445 69.110 63.815 69.120 ;
        RECT 63.445 68.850 64.465 69.110 ;
        RECT 67.615 68.930 68.255 69.140 ;
        RECT 63.445 68.840 63.815 68.850 ;
        RECT 66.550 68.810 68.255 68.930 ;
        RECT 68.770 69.110 69.140 69.120 ;
        RECT 68.770 68.850 69.790 69.110 ;
        RECT 72.940 68.930 73.580 69.140 ;
        RECT 78.275 68.930 78.915 69.140 ;
        RECT 68.770 68.840 69.140 68.850 ;
        RECT 71.875 68.810 73.580 68.930 ;
        RECT 77.210 68.810 78.915 68.930 ;
        RECT 79.430 69.110 79.800 69.120 ;
        RECT 79.430 68.850 80.450 69.110 ;
        RECT 83.600 68.930 84.240 69.140 ;
        RECT 79.430 68.840 79.800 68.850 ;
        RECT 82.535 68.810 84.240 68.930 ;
        RECT 84.765 69.110 85.135 69.120 ;
        RECT 84.765 68.850 85.785 69.110 ;
        RECT 88.935 68.930 89.575 69.140 ;
        RECT 84.765 68.840 85.135 68.850 ;
        RECT 87.870 68.810 89.575 68.930 ;
        RECT 90.090 69.110 90.460 69.120 ;
        RECT 90.090 68.850 91.110 69.110 ;
        RECT 94.260 68.930 94.900 69.140 ;
        RECT 90.090 68.840 90.460 68.850 ;
        RECT 93.195 68.810 94.900 68.930 ;
        RECT 95.425 69.110 95.795 69.120 ;
        RECT 95.425 68.850 96.445 69.110 ;
        RECT 99.595 68.930 100.235 69.140 ;
        RECT 95.425 68.840 95.795 68.850 ;
        RECT 98.530 68.810 100.235 68.930 ;
        RECT 100.750 69.110 101.120 69.120 ;
        RECT 100.750 68.850 101.770 69.110 ;
        RECT 104.920 68.930 105.560 69.140 ;
        RECT 100.750 68.840 101.120 68.850 ;
        RECT 103.855 68.810 105.560 68.930 ;
        RECT 106.085 69.110 106.455 69.120 ;
        RECT 106.085 68.850 107.105 69.110 ;
        RECT 110.255 68.930 110.895 69.140 ;
        RECT 106.085 68.840 106.455 68.850 ;
        RECT 109.190 68.810 110.895 68.930 ;
        RECT 111.410 69.110 111.780 69.120 ;
        RECT 111.410 68.850 112.430 69.110 ;
        RECT 115.580 68.930 116.220 69.140 ;
        RECT 120.915 68.930 121.555 69.140 ;
        RECT 111.410 68.840 111.780 68.850 ;
        RECT 114.515 68.810 116.220 68.930 ;
        RECT 119.850 68.810 121.555 68.930 ;
        RECT 38.095 68.670 41.600 68.810 ;
        RECT 43.430 68.670 46.935 68.810 ;
        RECT 48.755 68.670 52.260 68.810 ;
        RECT 54.090 68.670 57.595 68.810 ;
        RECT 59.415 68.670 62.920 68.810 ;
        RECT 64.750 68.670 68.255 68.810 ;
        RECT 70.075 68.670 73.580 68.810 ;
        RECT 75.410 68.670 78.915 68.810 ;
        RECT 80.735 68.670 84.240 68.810 ;
        RECT 86.070 68.670 89.575 68.810 ;
        RECT 91.395 68.670 94.900 68.810 ;
        RECT 96.730 68.670 100.235 68.810 ;
        RECT 102.055 68.670 105.560 68.810 ;
        RECT 107.390 68.670 110.895 68.810 ;
        RECT 112.715 68.670 116.220 68.810 ;
        RECT 118.050 68.670 121.555 68.810 ;
        RECT 36.840 68.350 41.600 68.670 ;
        RECT 42.175 68.350 46.935 68.670 ;
        RECT 47.500 68.350 52.260 68.670 ;
        RECT 52.835 68.350 57.595 68.670 ;
        RECT 58.160 68.350 62.920 68.670 ;
        RECT 63.495 68.350 68.255 68.670 ;
        RECT 68.820 68.350 73.580 68.670 ;
        RECT 74.155 68.350 78.915 68.670 ;
        RECT 79.480 68.350 84.240 68.670 ;
        RECT 84.815 68.350 89.575 68.670 ;
        RECT 90.140 68.350 94.900 68.670 ;
        RECT 95.475 68.350 100.235 68.670 ;
        RECT 100.800 68.350 105.560 68.670 ;
        RECT 106.135 68.350 110.895 68.670 ;
        RECT 111.460 68.350 116.220 68.670 ;
        RECT 116.795 68.350 121.555 68.670 ;
        RECT 32.040 68.000 34.915 68.260 ;
        RECT 32.040 67.830 32.300 68.000 ;
        RECT 31.480 67.570 32.300 67.830 ;
        RECT 34.655 67.825 34.915 68.000 ;
        RECT 36.840 68.210 40.345 68.350 ;
        RECT 42.175 68.210 45.680 68.350 ;
        RECT 47.500 68.210 51.005 68.350 ;
        RECT 52.835 68.210 56.340 68.350 ;
        RECT 58.160 68.210 61.665 68.350 ;
        RECT 63.495 68.210 67.000 68.350 ;
        RECT 68.820 68.210 72.325 68.350 ;
        RECT 74.155 68.210 77.660 68.350 ;
        RECT 79.480 68.210 82.985 68.350 ;
        RECT 84.815 68.210 88.320 68.350 ;
        RECT 90.140 68.210 93.645 68.350 ;
        RECT 95.475 68.210 98.980 68.350 ;
        RECT 100.800 68.210 104.305 68.350 ;
        RECT 106.135 68.210 109.640 68.350 ;
        RECT 111.460 68.210 114.965 68.350 ;
        RECT 116.795 68.210 120.300 68.350 ;
        RECT 36.840 68.090 38.545 68.210 ;
        RECT 41.285 68.160 41.655 68.170 ;
        RECT 32.625 67.485 34.390 67.765 ;
        RECT 34.655 67.565 36.305 67.825 ;
        RECT 36.840 67.615 37.480 68.090 ;
        RECT 40.580 67.900 41.655 68.160 ;
        RECT 41.285 67.890 41.655 67.900 ;
        RECT 42.175 68.090 43.880 68.210 ;
        RECT 46.620 68.160 46.990 68.170 ;
        RECT 37.950 67.485 38.320 67.765 ;
        RECT 38.715 67.485 39.110 67.765 ;
        RECT 39.330 67.485 39.730 67.765 ;
        RECT 42.175 67.615 42.815 68.090 ;
        RECT 45.915 67.900 46.990 68.160 ;
        RECT 46.620 67.890 46.990 67.900 ;
        RECT 47.500 68.090 49.205 68.210 ;
        RECT 51.945 68.160 52.315 68.170 ;
        RECT 43.285 67.485 43.655 67.765 ;
        RECT 44.050 67.485 44.445 67.765 ;
        RECT 44.665 67.485 45.065 67.765 ;
        RECT 47.500 67.615 48.140 68.090 ;
        RECT 51.240 67.900 52.315 68.160 ;
        RECT 51.945 67.890 52.315 67.900 ;
        RECT 52.835 68.090 54.540 68.210 ;
        RECT 57.280 68.160 57.650 68.170 ;
        RECT 48.610 67.485 48.980 67.765 ;
        RECT 49.375 67.485 49.770 67.765 ;
        RECT 49.990 67.485 50.390 67.765 ;
        RECT 52.835 67.615 53.475 68.090 ;
        RECT 56.575 67.900 57.650 68.160 ;
        RECT 57.280 67.890 57.650 67.900 ;
        RECT 58.160 68.090 59.865 68.210 ;
        RECT 62.605 68.160 62.975 68.170 ;
        RECT 54.710 67.485 55.105 67.765 ;
        RECT 55.325 67.485 55.725 67.765 ;
        RECT 58.160 67.615 58.800 68.090 ;
        RECT 61.900 67.900 62.975 68.160 ;
        RECT 62.605 67.890 62.975 67.900 ;
        RECT 63.495 68.090 65.200 68.210 ;
        RECT 67.940 68.160 68.310 68.170 ;
        RECT 59.270 67.485 59.640 67.765 ;
        RECT 60.035 67.485 60.430 67.765 ;
        RECT 60.650 67.485 61.050 67.765 ;
        RECT 63.495 67.615 64.135 68.090 ;
        RECT 67.235 67.900 68.310 68.160 ;
        RECT 67.940 67.890 68.310 67.900 ;
        RECT 68.820 68.090 70.525 68.210 ;
        RECT 73.265 68.160 73.635 68.170 ;
        RECT 64.605 67.485 64.975 67.765 ;
        RECT 65.370 67.485 65.765 67.765 ;
        RECT 65.985 67.485 66.385 67.765 ;
        RECT 68.820 67.615 69.460 68.090 ;
        RECT 72.560 67.900 73.635 68.160 ;
        RECT 73.265 67.890 73.635 67.900 ;
        RECT 74.155 68.090 75.860 68.210 ;
        RECT 78.600 68.160 78.970 68.170 ;
        RECT 69.930 67.485 70.300 67.765 ;
        RECT 70.695 67.485 71.090 67.765 ;
        RECT 71.310 67.485 71.710 67.765 ;
        RECT 74.155 67.615 74.795 68.090 ;
        RECT 77.895 67.900 78.970 68.160 ;
        RECT 78.600 67.890 78.970 67.900 ;
        RECT 79.480 68.090 81.185 68.210 ;
        RECT 83.925 68.160 84.295 68.170 ;
        RECT 75.265 67.485 76.425 67.765 ;
        RECT 76.645 67.485 77.045 67.765 ;
        RECT 79.480 67.615 80.120 68.090 ;
        RECT 83.220 67.900 84.295 68.160 ;
        RECT 83.925 67.890 84.295 67.900 ;
        RECT 84.815 68.090 86.520 68.210 ;
        RECT 89.260 68.160 89.630 68.170 ;
        RECT 80.590 67.485 80.960 67.765 ;
        RECT 81.355 67.485 81.750 67.765 ;
        RECT 81.970 67.485 82.370 67.765 ;
        RECT 84.815 67.615 85.455 68.090 ;
        RECT 88.555 67.900 89.630 68.160 ;
        RECT 89.260 67.890 89.630 67.900 ;
        RECT 90.140 68.090 91.845 68.210 ;
        RECT 94.585 68.160 94.955 68.170 ;
        RECT 85.925 67.485 86.295 67.765 ;
        RECT 86.690 67.485 87.085 67.765 ;
        RECT 87.305 67.485 87.705 67.765 ;
        RECT 90.140 67.615 90.780 68.090 ;
        RECT 93.880 67.900 94.955 68.160 ;
        RECT 94.585 67.890 94.955 67.900 ;
        RECT 95.475 68.090 97.180 68.210 ;
        RECT 99.920 68.160 100.290 68.170 ;
        RECT 91.250 67.485 91.620 67.765 ;
        RECT 92.015 67.485 92.410 67.765 ;
        RECT 92.630 67.485 93.030 67.765 ;
        RECT 95.475 67.615 96.115 68.090 ;
        RECT 99.215 67.900 100.290 68.160 ;
        RECT 99.920 67.890 100.290 67.900 ;
        RECT 100.800 68.090 102.505 68.210 ;
        RECT 105.245 68.160 105.615 68.170 ;
        RECT 97.350 67.485 97.745 67.765 ;
        RECT 97.965 67.485 98.365 67.765 ;
        RECT 100.800 67.615 101.440 68.090 ;
        RECT 104.540 67.900 105.615 68.160 ;
        RECT 105.245 67.890 105.615 67.900 ;
        RECT 106.135 68.090 107.840 68.210 ;
        RECT 110.580 68.160 110.950 68.170 ;
        RECT 101.910 67.485 102.280 67.765 ;
        RECT 102.675 67.485 103.070 67.765 ;
        RECT 103.290 67.485 103.690 67.765 ;
        RECT 106.135 67.615 106.775 68.090 ;
        RECT 109.875 67.900 110.950 68.160 ;
        RECT 110.580 67.890 110.950 67.900 ;
        RECT 111.460 68.090 113.165 68.210 ;
        RECT 115.905 68.160 116.275 68.170 ;
        RECT 107.245 67.485 107.615 67.765 ;
        RECT 108.010 67.485 108.405 67.765 ;
        RECT 108.625 67.485 109.025 67.765 ;
        RECT 111.460 67.615 112.100 68.090 ;
        RECT 115.200 67.900 116.275 68.160 ;
        RECT 115.905 67.890 116.275 67.900 ;
        RECT 116.795 68.090 118.500 68.210 ;
        RECT 121.240 68.160 121.610 68.170 ;
        RECT 112.570 67.485 112.940 67.765 ;
        RECT 113.335 67.485 113.730 67.765 ;
        RECT 113.950 67.485 114.350 67.765 ;
        RECT 116.795 67.615 117.435 68.090 ;
        RECT 120.535 67.900 121.610 68.160 ;
        RECT 121.240 67.890 121.610 67.900 ;
        RECT 122.645 68.000 125.520 68.260 ;
        RECT 122.645 67.830 122.905 68.000 ;
        RECT 117.905 67.485 119.065 67.765 ;
        RECT 119.285 67.485 119.685 67.765 ;
        RECT 122.085 67.570 122.905 67.830 ;
        RECT 125.260 67.825 125.520 68.000 ;
        RECT 123.230 67.485 124.995 67.765 ;
        RECT 125.260 67.565 126.910 67.825 ;
        RECT 36.785 67.265 37.155 67.275 ;
        RECT 42.120 67.265 42.490 67.275 ;
        RECT 47.445 67.265 47.815 67.275 ;
        RECT 52.780 67.265 53.150 67.275 ;
        RECT 58.105 67.265 58.475 67.275 ;
        RECT 63.440 67.265 63.810 67.275 ;
        RECT 68.765 67.265 69.135 67.275 ;
        RECT 79.425 67.265 79.795 67.275 ;
        RECT 84.760 67.265 85.130 67.275 ;
        RECT 90.085 67.265 90.455 67.275 ;
        RECT 95.420 67.265 95.790 67.275 ;
        RECT 100.745 67.265 101.115 67.275 ;
        RECT 106.080 67.265 106.450 67.275 ;
        RECT 111.405 67.265 111.775 67.275 ;
        RECT 36.785 67.005 37.810 67.265 ;
        RECT 41.285 67.175 41.655 67.185 ;
        RECT 36.785 66.995 37.155 67.005 ;
        RECT 28.415 66.555 28.695 66.925 ;
        RECT 40.630 66.915 41.655 67.175 ;
        RECT 42.120 67.005 43.145 67.265 ;
        RECT 46.620 67.175 46.990 67.185 ;
        RECT 42.120 66.995 42.490 67.005 ;
        RECT 45.965 66.915 46.990 67.175 ;
        RECT 47.445 67.005 48.470 67.265 ;
        RECT 51.945 67.175 52.315 67.185 ;
        RECT 47.445 66.995 47.815 67.005 ;
        RECT 51.290 66.915 52.315 67.175 ;
        RECT 52.780 67.005 53.805 67.265 ;
        RECT 57.280 67.175 57.650 67.185 ;
        RECT 52.780 66.995 53.150 67.005 ;
        RECT 56.625 66.915 57.650 67.175 ;
        RECT 58.105 67.005 59.130 67.265 ;
        RECT 62.605 67.175 62.975 67.185 ;
        RECT 58.105 66.995 58.475 67.005 ;
        RECT 61.950 66.915 62.975 67.175 ;
        RECT 63.440 67.005 64.465 67.265 ;
        RECT 67.940 67.175 68.310 67.185 ;
        RECT 63.440 66.995 63.810 67.005 ;
        RECT 67.285 66.915 68.310 67.175 ;
        RECT 68.765 67.005 69.790 67.265 ;
        RECT 73.265 67.175 73.635 67.185 ;
        RECT 78.600 67.175 78.970 67.185 ;
        RECT 68.765 66.995 69.135 67.005 ;
        RECT 72.610 66.915 73.635 67.175 ;
        RECT 77.945 66.915 78.970 67.175 ;
        RECT 79.425 67.005 80.450 67.265 ;
        RECT 83.925 67.175 84.295 67.185 ;
        RECT 79.425 66.995 79.795 67.005 ;
        RECT 83.270 66.915 84.295 67.175 ;
        RECT 84.760 67.005 85.785 67.265 ;
        RECT 89.260 67.175 89.630 67.185 ;
        RECT 84.760 66.995 85.130 67.005 ;
        RECT 88.605 66.915 89.630 67.175 ;
        RECT 90.085 67.005 91.110 67.265 ;
        RECT 94.585 67.175 94.955 67.185 ;
        RECT 90.085 66.995 90.455 67.005 ;
        RECT 93.930 66.915 94.955 67.175 ;
        RECT 95.420 67.005 96.445 67.265 ;
        RECT 99.920 67.175 100.290 67.185 ;
        RECT 95.420 66.995 95.790 67.005 ;
        RECT 99.265 66.915 100.290 67.175 ;
        RECT 100.745 67.005 101.770 67.265 ;
        RECT 105.245 67.175 105.615 67.185 ;
        RECT 100.745 66.995 101.115 67.005 ;
        RECT 104.590 66.915 105.615 67.175 ;
        RECT 106.080 67.005 107.105 67.265 ;
        RECT 110.580 67.175 110.950 67.185 ;
        RECT 106.080 66.995 106.450 67.005 ;
        RECT 109.925 66.915 110.950 67.175 ;
        RECT 111.405 67.005 112.430 67.265 ;
        RECT 115.905 67.175 116.275 67.185 ;
        RECT 121.240 67.175 121.610 67.185 ;
        RECT 111.405 66.995 111.775 67.005 ;
        RECT 115.250 66.915 116.275 67.175 ;
        RECT 120.585 66.915 121.610 67.175 ;
        RECT 41.285 66.905 41.655 66.915 ;
        RECT 46.620 66.905 46.990 66.915 ;
        RECT 51.945 66.905 52.315 66.915 ;
        RECT 57.280 66.905 57.650 66.915 ;
        RECT 62.605 66.905 62.975 66.915 ;
        RECT 67.940 66.905 68.310 66.915 ;
        RECT 73.265 66.905 73.635 66.915 ;
        RECT 78.600 66.905 78.970 66.915 ;
        RECT 83.925 66.905 84.295 66.915 ;
        RECT 89.260 66.905 89.630 66.915 ;
        RECT 94.585 66.905 94.955 66.915 ;
        RECT 99.920 66.905 100.290 66.915 ;
        RECT 105.245 66.905 105.615 66.915 ;
        RECT 110.580 66.905 110.950 66.915 ;
        RECT 115.905 66.905 116.275 66.915 ;
        RECT 121.240 66.905 121.610 66.915 ;
        RECT 28.030 65.225 28.310 65.595 ;
        RECT 27.655 63.285 27.935 63.655 ;
        RECT 27.270 60.955 27.550 61.325 ;
        RECT 26.895 55.750 27.175 56.120 ;
        RECT 26.510 53.420 26.790 53.790 ;
        RECT 26.135 41.970 26.415 42.340 ;
        RECT 25.755 40.680 26.035 41.050 ;
        RECT 25.385 39.185 25.645 40.295 ;
        RECT 14.605 35.880 15.985 36.170 ;
        RECT 25.005 35.465 25.265 36.570 ;
        RECT 10.530 27.500 10.790 33.015 ;
        RECT 11.745 32.495 13.345 32.785 ;
        RECT 12.430 26.945 12.690 32.495 ;
        RECT 16.040 32.050 17.645 32.340 ;
        RECT 16.110 31.490 16.565 32.050 ;
        RECT 15.455 31.035 16.565 31.490 ;
        RECT 15.455 28.030 15.910 31.035 ;
        RECT 14.605 27.740 15.985 28.030 ;
        RECT 10.530 19.360 10.790 24.875 ;
        RECT 11.745 24.355 13.345 24.645 ;
        RECT 12.430 18.805 12.690 24.355 ;
        RECT 16.040 23.910 17.645 24.200 ;
        RECT 16.110 23.350 16.565 23.910 ;
        RECT 15.455 22.895 16.565 23.350 ;
        RECT 15.455 19.890 15.910 22.895 ;
        RECT 14.605 19.600 15.985 19.890 ;
        RECT 10.530 11.220 10.790 16.735 ;
        RECT 11.745 16.215 13.345 16.505 ;
        RECT 12.430 10.665 12.690 16.215 ;
        RECT 16.040 15.770 17.645 16.060 ;
        RECT 16.110 15.210 16.565 15.770 ;
        RECT 15.455 14.755 16.565 15.210 ;
        RECT 15.455 11.750 15.910 14.755 ;
        RECT 25.045 12.200 25.225 35.465 ;
        RECT 24.995 11.830 25.275 12.200 ;
        RECT 14.605 11.460 15.985 11.750 ;
        RECT 25.425 10.910 25.605 39.185 ;
        RECT 25.805 37.430 25.985 40.680 ;
        RECT 26.185 38.720 26.365 41.970 ;
        RECT 26.130 38.350 26.410 38.720 ;
        RECT 25.755 37.060 26.035 37.430 ;
        RECT 25.805 28.430 25.985 37.060 ;
        RECT 26.185 33.155 26.365 38.350 ;
        RECT 26.145 32.045 26.405 33.155 ;
        RECT 26.185 32.000 26.365 32.045 ;
        RECT 25.765 27.325 26.025 28.430 ;
        RECT 25.805 27.290 25.985 27.325 ;
        RECT 26.565 25.980 26.745 53.420 ;
        RECT 26.945 52.500 27.125 55.750 ;
        RECT 26.895 52.130 27.175 52.500 ;
        RECT 26.945 27.270 27.125 52.130 ;
        RECT 27.325 48.585 27.505 60.955 ;
        RECT 27.705 60.035 27.885 63.285 ;
        RECT 27.655 59.665 27.935 60.035 ;
        RECT 27.705 49.875 27.885 59.665 ;
        RECT 28.085 59.390 28.265 65.225 ;
        RECT 28.465 64.300 28.645 66.555 ;
        RECT 36.785 65.240 37.155 65.250 ;
        RECT 42.120 65.240 42.490 65.250 ;
        RECT 47.445 65.240 47.815 65.250 ;
        RECT 52.780 65.240 53.150 65.250 ;
        RECT 58.105 65.240 58.475 65.250 ;
        RECT 63.440 65.240 63.810 65.250 ;
        RECT 68.765 65.240 69.135 65.250 ;
        RECT 74.100 65.240 74.470 65.250 ;
        RECT 79.425 65.240 79.795 65.250 ;
        RECT 84.760 65.240 85.130 65.250 ;
        RECT 90.085 65.240 90.455 65.250 ;
        RECT 95.420 65.240 95.790 65.250 ;
        RECT 100.745 65.240 101.115 65.250 ;
        RECT 106.080 65.240 106.450 65.250 ;
        RECT 111.405 65.240 111.775 65.250 ;
        RECT 116.740 65.240 117.110 65.250 ;
        RECT 36.785 64.980 37.810 65.240 ;
        RECT 41.285 65.145 41.655 65.155 ;
        RECT 36.785 64.970 37.155 64.980 ;
        RECT 40.630 64.885 41.655 65.145 ;
        RECT 42.120 64.980 43.145 65.240 ;
        RECT 46.620 65.145 46.990 65.155 ;
        RECT 42.120 64.970 42.490 64.980 ;
        RECT 45.965 64.885 46.990 65.145 ;
        RECT 47.445 64.980 48.470 65.240 ;
        RECT 51.945 65.145 52.315 65.155 ;
        RECT 47.445 64.970 47.815 64.980 ;
        RECT 51.290 64.885 52.315 65.145 ;
        RECT 52.780 64.980 53.805 65.240 ;
        RECT 57.280 65.145 57.650 65.155 ;
        RECT 52.780 64.970 53.150 64.980 ;
        RECT 56.625 64.885 57.650 65.145 ;
        RECT 58.105 64.980 59.130 65.240 ;
        RECT 62.605 65.145 62.975 65.155 ;
        RECT 58.105 64.970 58.475 64.980 ;
        RECT 61.950 64.885 62.975 65.145 ;
        RECT 63.440 64.980 64.465 65.240 ;
        RECT 67.940 65.145 68.310 65.155 ;
        RECT 63.440 64.970 63.810 64.980 ;
        RECT 67.285 64.885 68.310 65.145 ;
        RECT 68.765 64.980 69.790 65.240 ;
        RECT 73.265 65.145 73.635 65.155 ;
        RECT 68.765 64.970 69.135 64.980 ;
        RECT 72.610 64.885 73.635 65.145 ;
        RECT 74.100 64.980 75.125 65.240 ;
        RECT 78.600 65.145 78.970 65.155 ;
        RECT 74.100 64.970 74.470 64.980 ;
        RECT 77.945 64.885 78.970 65.145 ;
        RECT 79.425 64.980 80.450 65.240 ;
        RECT 83.925 65.145 84.295 65.155 ;
        RECT 79.425 64.970 79.795 64.980 ;
        RECT 83.270 64.885 84.295 65.145 ;
        RECT 84.760 64.980 85.785 65.240 ;
        RECT 89.260 65.145 89.630 65.155 ;
        RECT 84.760 64.970 85.130 64.980 ;
        RECT 88.605 64.885 89.630 65.145 ;
        RECT 90.085 64.980 91.110 65.240 ;
        RECT 94.585 65.145 94.955 65.155 ;
        RECT 90.085 64.970 90.455 64.980 ;
        RECT 93.930 64.885 94.955 65.145 ;
        RECT 95.420 64.980 96.445 65.240 ;
        RECT 99.920 65.145 100.290 65.155 ;
        RECT 95.420 64.970 95.790 64.980 ;
        RECT 99.265 64.885 100.290 65.145 ;
        RECT 100.745 64.980 101.770 65.240 ;
        RECT 105.245 65.145 105.615 65.155 ;
        RECT 100.745 64.970 101.115 64.980 ;
        RECT 104.590 64.885 105.615 65.145 ;
        RECT 106.080 64.980 107.105 65.240 ;
        RECT 110.580 65.145 110.950 65.155 ;
        RECT 106.080 64.970 106.450 64.980 ;
        RECT 109.925 64.885 110.950 65.145 ;
        RECT 111.405 64.980 112.430 65.240 ;
        RECT 115.905 65.145 116.275 65.155 ;
        RECT 111.405 64.970 111.775 64.980 ;
        RECT 115.250 64.885 116.275 65.145 ;
        RECT 116.740 64.980 117.765 65.240 ;
        RECT 121.240 65.145 121.610 65.155 ;
        RECT 116.740 64.970 117.110 64.980 ;
        RECT 120.585 64.885 121.610 65.145 ;
        RECT 41.285 64.875 41.655 64.885 ;
        RECT 46.620 64.875 46.990 64.885 ;
        RECT 51.945 64.875 52.315 64.885 ;
        RECT 57.280 64.875 57.650 64.885 ;
        RECT 62.605 64.875 62.975 64.885 ;
        RECT 67.940 64.875 68.310 64.885 ;
        RECT 73.265 64.875 73.635 64.885 ;
        RECT 78.600 64.875 78.970 64.885 ;
        RECT 83.925 64.875 84.295 64.885 ;
        RECT 89.260 64.875 89.630 64.885 ;
        RECT 94.585 64.875 94.955 64.885 ;
        RECT 99.920 64.875 100.290 64.885 ;
        RECT 105.245 64.875 105.615 64.885 ;
        RECT 110.580 64.875 110.950 64.885 ;
        RECT 115.905 64.875 116.275 64.885 ;
        RECT 121.240 64.875 121.610 64.885 ;
        RECT 34.005 64.590 34.400 64.595 ;
        RECT 33.390 64.310 35.160 64.590 ;
        RECT 38.715 64.310 39.110 64.590 ;
        RECT 39.330 64.315 39.730 64.595 ;
        RECT 40.015 64.310 40.485 64.590 ;
        RECT 44.050 64.310 44.445 64.590 ;
        RECT 44.665 64.315 45.065 64.595 ;
        RECT 45.350 64.310 45.820 64.590 ;
        RECT 49.375 64.310 49.770 64.590 ;
        RECT 49.990 64.315 50.390 64.595 ;
        RECT 50.675 64.310 51.145 64.590 ;
        RECT 54.710 64.310 55.105 64.590 ;
        RECT 55.325 64.315 55.725 64.595 ;
        RECT 56.010 64.310 56.480 64.590 ;
        RECT 60.035 64.310 60.430 64.590 ;
        RECT 60.650 64.315 61.050 64.595 ;
        RECT 61.335 64.310 61.805 64.590 ;
        RECT 65.370 64.310 65.765 64.590 ;
        RECT 65.985 64.315 66.385 64.595 ;
        RECT 66.670 64.310 67.140 64.590 ;
        RECT 70.695 64.310 71.090 64.590 ;
        RECT 71.310 64.315 71.710 64.595 ;
        RECT 71.995 64.310 72.465 64.590 ;
        RECT 76.030 64.310 76.425 64.590 ;
        RECT 76.645 64.315 77.045 64.595 ;
        RECT 77.330 64.310 77.800 64.590 ;
        RECT 81.355 64.310 81.750 64.590 ;
        RECT 81.970 64.315 82.370 64.595 ;
        RECT 82.655 64.310 83.125 64.590 ;
        RECT 86.690 64.310 87.085 64.590 ;
        RECT 87.305 64.315 87.705 64.595 ;
        RECT 87.990 64.310 88.460 64.590 ;
        RECT 92.015 64.310 92.410 64.590 ;
        RECT 92.630 64.315 93.030 64.595 ;
        RECT 93.315 64.310 93.785 64.590 ;
        RECT 97.350 64.310 97.745 64.590 ;
        RECT 97.965 64.315 98.365 64.595 ;
        RECT 98.650 64.310 99.120 64.590 ;
        RECT 102.675 64.310 103.070 64.590 ;
        RECT 103.290 64.315 103.690 64.595 ;
        RECT 103.975 64.310 104.445 64.590 ;
        RECT 108.010 64.310 108.405 64.590 ;
        RECT 108.625 64.315 109.025 64.595 ;
        RECT 109.310 64.310 109.780 64.590 ;
        RECT 113.335 64.310 113.730 64.590 ;
        RECT 113.950 64.315 114.350 64.595 ;
        RECT 114.635 64.310 115.105 64.590 ;
        RECT 118.670 64.310 119.065 64.590 ;
        RECT 119.285 64.315 119.685 64.595 ;
        RECT 124.610 64.590 125.005 64.595 ;
        RECT 119.970 64.310 120.440 64.590 ;
        RECT 123.995 64.310 125.765 64.590 ;
        RECT 28.415 63.930 28.695 64.300 ;
        RECT 36.785 63.940 37.155 63.950 ;
        RECT 42.120 63.940 42.490 63.950 ;
        RECT 47.445 63.940 47.815 63.950 ;
        RECT 52.780 63.940 53.150 63.950 ;
        RECT 58.105 63.940 58.475 63.950 ;
        RECT 63.440 63.940 63.810 63.950 ;
        RECT 68.765 63.940 69.135 63.950 ;
        RECT 74.100 63.940 74.470 63.950 ;
        RECT 79.425 63.940 79.795 63.950 ;
        RECT 84.760 63.940 85.130 63.950 ;
        RECT 90.085 63.940 90.455 63.950 ;
        RECT 95.420 63.940 95.790 63.950 ;
        RECT 100.745 63.940 101.115 63.950 ;
        RECT 106.080 63.940 106.450 63.950 ;
        RECT 111.405 63.940 111.775 63.950 ;
        RECT 116.740 63.940 117.110 63.950 ;
        RECT 28.465 60.680 28.645 63.930 ;
        RECT 36.785 63.680 37.860 63.940 ;
        RECT 42.120 63.680 43.195 63.940 ;
        RECT 47.445 63.680 48.520 63.940 ;
        RECT 52.780 63.680 53.855 63.940 ;
        RECT 58.105 63.680 59.180 63.940 ;
        RECT 63.440 63.680 64.515 63.940 ;
        RECT 68.765 63.680 69.840 63.940 ;
        RECT 74.100 63.680 75.175 63.940 ;
        RECT 79.425 63.680 80.500 63.940 ;
        RECT 84.760 63.680 85.835 63.940 ;
        RECT 90.085 63.680 91.160 63.940 ;
        RECT 95.420 63.680 96.495 63.940 ;
        RECT 100.745 63.680 101.820 63.940 ;
        RECT 106.080 63.680 107.155 63.940 ;
        RECT 111.405 63.680 112.480 63.940 ;
        RECT 116.740 63.680 117.815 63.940 ;
        RECT 36.785 63.670 37.155 63.680 ;
        RECT 42.120 63.670 42.490 63.680 ;
        RECT 47.445 63.670 47.815 63.680 ;
        RECT 52.780 63.670 53.150 63.680 ;
        RECT 58.105 63.670 58.475 63.680 ;
        RECT 63.440 63.670 63.810 63.680 ;
        RECT 68.765 63.670 69.135 63.680 ;
        RECT 74.100 63.670 74.470 63.680 ;
        RECT 79.425 63.670 79.795 63.680 ;
        RECT 84.760 63.670 85.130 63.680 ;
        RECT 90.085 63.670 90.455 63.680 ;
        RECT 95.420 63.670 95.790 63.680 ;
        RECT 100.745 63.670 101.115 63.680 ;
        RECT 106.080 63.670 106.450 63.680 ;
        RECT 111.405 63.670 111.775 63.680 ;
        RECT 116.740 63.670 117.110 63.680 ;
        RECT 41.290 63.310 41.660 63.320 ;
        RECT 46.625 63.310 46.995 63.320 ;
        RECT 51.950 63.310 52.320 63.320 ;
        RECT 57.285 63.310 57.655 63.320 ;
        RECT 62.610 63.310 62.980 63.320 ;
        RECT 67.945 63.310 68.315 63.320 ;
        RECT 73.270 63.310 73.640 63.320 ;
        RECT 78.605 63.310 78.975 63.320 ;
        RECT 83.930 63.310 84.300 63.320 ;
        RECT 89.265 63.310 89.635 63.320 ;
        RECT 94.590 63.310 94.960 63.320 ;
        RECT 99.925 63.310 100.295 63.320 ;
        RECT 105.250 63.310 105.620 63.320 ;
        RECT 110.585 63.310 110.955 63.320 ;
        RECT 115.910 63.310 116.280 63.320 ;
        RECT 121.245 63.310 121.615 63.320 ;
        RECT 40.630 63.050 41.660 63.310 ;
        RECT 45.965 63.050 46.995 63.310 ;
        RECT 51.290 63.050 52.320 63.310 ;
        RECT 56.625 63.050 57.655 63.310 ;
        RECT 61.950 63.050 62.980 63.310 ;
        RECT 67.285 63.050 68.315 63.310 ;
        RECT 72.610 63.050 73.640 63.310 ;
        RECT 77.945 63.050 78.975 63.310 ;
        RECT 83.270 63.050 84.300 63.310 ;
        RECT 88.605 63.050 89.635 63.310 ;
        RECT 93.930 63.050 94.960 63.310 ;
        RECT 99.265 63.050 100.295 63.310 ;
        RECT 104.590 63.050 105.620 63.310 ;
        RECT 109.925 63.050 110.955 63.310 ;
        RECT 115.250 63.050 116.280 63.310 ;
        RECT 120.585 63.050 121.615 63.310 ;
        RECT 41.290 63.040 41.660 63.050 ;
        RECT 46.625 63.040 46.995 63.050 ;
        RECT 51.950 63.040 52.320 63.050 ;
        RECT 57.285 63.040 57.655 63.050 ;
        RECT 62.610 63.040 62.980 63.050 ;
        RECT 67.945 63.040 68.315 63.050 ;
        RECT 73.270 63.040 73.640 63.050 ;
        RECT 78.605 63.040 78.975 63.050 ;
        RECT 83.930 63.040 84.300 63.050 ;
        RECT 89.265 63.040 89.635 63.050 ;
        RECT 94.590 63.040 94.960 63.050 ;
        RECT 99.925 63.040 100.295 63.050 ;
        RECT 105.250 63.040 105.620 63.050 ;
        RECT 110.585 63.040 110.955 63.050 ;
        RECT 115.910 63.040 116.280 63.050 ;
        RECT 121.245 63.040 121.615 63.050 ;
        RECT 36.790 61.575 37.160 61.585 ;
        RECT 42.125 61.575 42.495 61.585 ;
        RECT 47.450 61.575 47.820 61.585 ;
        RECT 52.785 61.575 53.155 61.585 ;
        RECT 58.110 61.575 58.480 61.585 ;
        RECT 63.445 61.575 63.815 61.585 ;
        RECT 68.770 61.575 69.140 61.585 ;
        RECT 74.105 61.575 74.475 61.585 ;
        RECT 79.430 61.575 79.800 61.585 ;
        RECT 84.765 61.575 85.135 61.585 ;
        RECT 90.090 61.575 90.460 61.585 ;
        RECT 95.425 61.575 95.795 61.585 ;
        RECT 100.750 61.575 101.120 61.585 ;
        RECT 106.085 61.575 106.455 61.585 ;
        RECT 111.410 61.575 111.780 61.585 ;
        RECT 116.745 61.575 117.115 61.585 ;
        RECT 36.790 61.315 37.810 61.575 ;
        RECT 42.125 61.315 43.145 61.575 ;
        RECT 47.450 61.315 48.470 61.575 ;
        RECT 52.785 61.315 53.805 61.575 ;
        RECT 58.110 61.315 59.130 61.575 ;
        RECT 63.445 61.315 64.465 61.575 ;
        RECT 68.770 61.315 69.790 61.575 ;
        RECT 74.105 61.315 75.125 61.575 ;
        RECT 79.430 61.315 80.450 61.575 ;
        RECT 84.765 61.315 85.785 61.575 ;
        RECT 90.090 61.315 91.110 61.575 ;
        RECT 95.425 61.315 96.445 61.575 ;
        RECT 100.750 61.315 101.770 61.575 ;
        RECT 106.085 61.315 107.105 61.575 ;
        RECT 111.410 61.315 112.430 61.575 ;
        RECT 116.745 61.315 117.765 61.575 ;
        RECT 36.790 61.305 37.160 61.315 ;
        RECT 42.125 61.305 42.495 61.315 ;
        RECT 47.450 61.305 47.820 61.315 ;
        RECT 52.785 61.305 53.155 61.315 ;
        RECT 58.110 61.305 58.480 61.315 ;
        RECT 63.445 61.305 63.815 61.315 ;
        RECT 68.770 61.305 69.140 61.315 ;
        RECT 74.105 61.305 74.475 61.315 ;
        RECT 79.430 61.305 79.800 61.315 ;
        RECT 84.765 61.305 85.135 61.315 ;
        RECT 90.090 61.305 90.460 61.315 ;
        RECT 95.425 61.305 95.795 61.315 ;
        RECT 100.750 61.305 101.120 61.315 ;
        RECT 106.085 61.305 106.455 61.315 ;
        RECT 111.410 61.305 111.780 61.315 ;
        RECT 116.745 61.305 117.115 61.315 ;
        RECT 41.285 60.925 41.655 60.935 ;
        RECT 46.620 60.925 46.990 60.935 ;
        RECT 51.945 60.925 52.315 60.935 ;
        RECT 57.280 60.925 57.650 60.935 ;
        RECT 62.605 60.925 62.975 60.935 ;
        RECT 67.940 60.925 68.310 60.935 ;
        RECT 73.265 60.925 73.635 60.935 ;
        RECT 78.600 60.925 78.970 60.935 ;
        RECT 83.925 60.925 84.295 60.935 ;
        RECT 89.260 60.925 89.630 60.935 ;
        RECT 94.585 60.925 94.955 60.935 ;
        RECT 99.920 60.925 100.290 60.935 ;
        RECT 105.245 60.925 105.615 60.935 ;
        RECT 110.580 60.925 110.950 60.935 ;
        RECT 115.905 60.925 116.275 60.935 ;
        RECT 121.240 60.925 121.610 60.935 ;
        RECT 28.415 60.310 28.695 60.680 ;
        RECT 40.580 60.665 41.655 60.925 ;
        RECT 45.915 60.665 46.990 60.925 ;
        RECT 51.240 60.665 52.315 60.925 ;
        RECT 56.575 60.665 57.650 60.925 ;
        RECT 61.900 60.665 62.975 60.925 ;
        RECT 67.235 60.665 68.310 60.925 ;
        RECT 72.560 60.665 73.635 60.925 ;
        RECT 77.895 60.665 78.970 60.925 ;
        RECT 83.220 60.665 84.295 60.925 ;
        RECT 88.555 60.665 89.630 60.925 ;
        RECT 93.880 60.665 94.955 60.925 ;
        RECT 99.215 60.665 100.290 60.925 ;
        RECT 104.540 60.665 105.615 60.925 ;
        RECT 109.875 60.665 110.950 60.925 ;
        RECT 115.200 60.665 116.275 60.925 ;
        RECT 120.535 60.665 121.610 60.925 ;
        RECT 41.285 60.655 41.655 60.665 ;
        RECT 46.620 60.655 46.990 60.665 ;
        RECT 51.945 60.655 52.315 60.665 ;
        RECT 57.280 60.655 57.650 60.665 ;
        RECT 62.605 60.655 62.975 60.665 ;
        RECT 67.940 60.655 68.310 60.665 ;
        RECT 73.265 60.655 73.635 60.665 ;
        RECT 78.600 60.655 78.970 60.665 ;
        RECT 83.925 60.655 84.295 60.665 ;
        RECT 89.260 60.655 89.630 60.665 ;
        RECT 94.585 60.655 94.955 60.665 ;
        RECT 99.920 60.655 100.290 60.665 ;
        RECT 105.245 60.655 105.615 60.665 ;
        RECT 110.580 60.655 110.950 60.665 ;
        RECT 115.905 60.655 116.275 60.665 ;
        RECT 121.240 60.655 121.610 60.665 ;
        RECT 28.035 59.020 28.315 59.390 ;
        RECT 28.085 56.765 28.265 59.020 ;
        RECT 28.465 58.060 28.645 60.310 ;
        RECT 32.625 59.950 34.390 60.230 ;
        RECT 37.950 59.950 38.470 60.230 ;
        RECT 38.715 59.950 39.110 60.230 ;
        RECT 39.330 59.950 39.730 60.230 ;
        RECT 43.285 59.950 43.805 60.230 ;
        RECT 44.050 59.950 44.445 60.230 ;
        RECT 44.665 59.950 45.065 60.230 ;
        RECT 48.610 59.950 49.130 60.230 ;
        RECT 49.375 59.950 49.770 60.230 ;
        RECT 49.990 59.950 50.390 60.230 ;
        RECT 53.945 59.950 54.465 60.230 ;
        RECT 54.710 59.950 55.105 60.230 ;
        RECT 55.325 59.950 55.725 60.230 ;
        RECT 59.270 59.950 59.790 60.230 ;
        RECT 60.035 59.950 60.430 60.230 ;
        RECT 60.650 59.950 61.050 60.230 ;
        RECT 64.605 59.950 65.125 60.230 ;
        RECT 65.370 59.950 65.765 60.230 ;
        RECT 65.985 59.950 66.385 60.230 ;
        RECT 69.930 59.950 70.450 60.230 ;
        RECT 70.695 59.950 71.090 60.230 ;
        RECT 71.310 59.950 71.710 60.230 ;
        RECT 75.265 59.950 75.785 60.230 ;
        RECT 76.030 59.950 76.425 60.230 ;
        RECT 76.645 59.950 77.045 60.230 ;
        RECT 80.590 59.950 81.110 60.230 ;
        RECT 81.355 59.950 81.750 60.230 ;
        RECT 81.970 59.950 82.370 60.230 ;
        RECT 85.925 59.950 86.445 60.230 ;
        RECT 86.690 59.950 87.085 60.230 ;
        RECT 87.305 59.950 87.705 60.230 ;
        RECT 91.250 59.950 91.770 60.230 ;
        RECT 92.015 59.950 92.410 60.230 ;
        RECT 92.630 59.950 93.030 60.230 ;
        RECT 96.585 59.950 97.105 60.230 ;
        RECT 97.350 59.950 97.745 60.230 ;
        RECT 97.965 59.950 98.365 60.230 ;
        RECT 101.910 59.950 102.430 60.230 ;
        RECT 102.675 59.950 103.070 60.230 ;
        RECT 103.290 59.950 103.690 60.230 ;
        RECT 107.245 59.950 107.765 60.230 ;
        RECT 108.010 59.950 108.405 60.230 ;
        RECT 108.625 59.950 109.025 60.230 ;
        RECT 112.570 59.950 113.090 60.230 ;
        RECT 113.335 59.950 113.730 60.230 ;
        RECT 113.950 59.950 114.350 60.230 ;
        RECT 117.905 59.950 118.425 60.230 ;
        RECT 118.670 59.950 119.065 60.230 ;
        RECT 119.285 59.950 119.685 60.230 ;
        RECT 123.230 59.950 124.995 60.230 ;
        RECT 36.785 59.730 37.155 59.740 ;
        RECT 42.120 59.730 42.490 59.740 ;
        RECT 47.445 59.730 47.815 59.740 ;
        RECT 52.780 59.730 53.150 59.740 ;
        RECT 58.105 59.730 58.475 59.740 ;
        RECT 63.440 59.730 63.810 59.740 ;
        RECT 68.765 59.730 69.135 59.740 ;
        RECT 74.100 59.730 74.470 59.740 ;
        RECT 79.425 59.730 79.795 59.740 ;
        RECT 84.760 59.730 85.130 59.740 ;
        RECT 90.085 59.730 90.455 59.740 ;
        RECT 95.420 59.730 95.790 59.740 ;
        RECT 100.745 59.730 101.115 59.740 ;
        RECT 106.080 59.730 106.450 59.740 ;
        RECT 111.405 59.730 111.775 59.740 ;
        RECT 116.740 59.730 117.110 59.740 ;
        RECT 36.785 59.470 37.810 59.730 ;
        RECT 41.285 59.640 41.655 59.650 ;
        RECT 36.785 59.460 37.155 59.470 ;
        RECT 40.630 59.380 41.655 59.640 ;
        RECT 42.120 59.470 43.145 59.730 ;
        RECT 46.620 59.640 46.990 59.650 ;
        RECT 42.120 59.460 42.490 59.470 ;
        RECT 45.965 59.380 46.990 59.640 ;
        RECT 47.445 59.470 48.470 59.730 ;
        RECT 51.945 59.640 52.315 59.650 ;
        RECT 47.445 59.460 47.815 59.470 ;
        RECT 51.290 59.380 52.315 59.640 ;
        RECT 52.780 59.470 53.805 59.730 ;
        RECT 57.280 59.640 57.650 59.650 ;
        RECT 52.780 59.460 53.150 59.470 ;
        RECT 56.625 59.380 57.650 59.640 ;
        RECT 58.105 59.470 59.130 59.730 ;
        RECT 62.605 59.640 62.975 59.650 ;
        RECT 58.105 59.460 58.475 59.470 ;
        RECT 61.950 59.380 62.975 59.640 ;
        RECT 63.440 59.470 64.465 59.730 ;
        RECT 67.940 59.640 68.310 59.650 ;
        RECT 63.440 59.460 63.810 59.470 ;
        RECT 67.285 59.380 68.310 59.640 ;
        RECT 68.765 59.470 69.790 59.730 ;
        RECT 73.265 59.640 73.635 59.650 ;
        RECT 68.765 59.460 69.135 59.470 ;
        RECT 72.610 59.380 73.635 59.640 ;
        RECT 74.100 59.470 75.125 59.730 ;
        RECT 78.600 59.640 78.970 59.650 ;
        RECT 74.100 59.460 74.470 59.470 ;
        RECT 77.945 59.380 78.970 59.640 ;
        RECT 79.425 59.470 80.450 59.730 ;
        RECT 83.925 59.640 84.295 59.650 ;
        RECT 79.425 59.460 79.795 59.470 ;
        RECT 83.270 59.380 84.295 59.640 ;
        RECT 84.760 59.470 85.785 59.730 ;
        RECT 89.260 59.640 89.630 59.650 ;
        RECT 84.760 59.460 85.130 59.470 ;
        RECT 88.605 59.380 89.630 59.640 ;
        RECT 90.085 59.470 91.110 59.730 ;
        RECT 94.585 59.640 94.955 59.650 ;
        RECT 90.085 59.460 90.455 59.470 ;
        RECT 93.930 59.380 94.955 59.640 ;
        RECT 95.420 59.470 96.445 59.730 ;
        RECT 99.920 59.640 100.290 59.650 ;
        RECT 95.420 59.460 95.790 59.470 ;
        RECT 99.265 59.380 100.290 59.640 ;
        RECT 100.745 59.470 101.770 59.730 ;
        RECT 105.245 59.640 105.615 59.650 ;
        RECT 100.745 59.460 101.115 59.470 ;
        RECT 104.590 59.380 105.615 59.640 ;
        RECT 106.080 59.470 107.105 59.730 ;
        RECT 110.580 59.640 110.950 59.650 ;
        RECT 106.080 59.460 106.450 59.470 ;
        RECT 109.925 59.380 110.950 59.640 ;
        RECT 111.405 59.470 112.430 59.730 ;
        RECT 115.905 59.640 116.275 59.650 ;
        RECT 111.405 59.460 111.775 59.470 ;
        RECT 115.250 59.380 116.275 59.640 ;
        RECT 116.740 59.470 117.765 59.730 ;
        RECT 121.240 59.640 121.610 59.650 ;
        RECT 116.740 59.460 117.110 59.470 ;
        RECT 120.585 59.380 121.610 59.640 ;
        RECT 41.285 59.370 41.655 59.380 ;
        RECT 46.620 59.370 46.990 59.380 ;
        RECT 51.945 59.370 52.315 59.380 ;
        RECT 57.280 59.370 57.650 59.380 ;
        RECT 62.605 59.370 62.975 59.380 ;
        RECT 67.940 59.370 68.310 59.380 ;
        RECT 73.265 59.370 73.635 59.380 ;
        RECT 78.600 59.370 78.970 59.380 ;
        RECT 83.925 59.370 84.295 59.380 ;
        RECT 89.260 59.370 89.630 59.380 ;
        RECT 94.585 59.370 94.955 59.380 ;
        RECT 99.920 59.370 100.290 59.380 ;
        RECT 105.245 59.370 105.615 59.380 ;
        RECT 110.580 59.370 110.950 59.380 ;
        RECT 115.905 59.370 116.275 59.380 ;
        RECT 121.240 59.370 121.610 59.380 ;
        RECT 28.410 57.690 28.690 58.060 ;
        RECT 36.785 57.705 37.155 57.715 ;
        RECT 42.120 57.705 42.490 57.715 ;
        RECT 47.445 57.705 47.815 57.715 ;
        RECT 52.780 57.705 53.150 57.715 ;
        RECT 58.105 57.705 58.475 57.715 ;
        RECT 63.440 57.705 63.810 57.715 ;
        RECT 68.765 57.705 69.135 57.715 ;
        RECT 74.100 57.705 74.470 57.715 ;
        RECT 79.425 57.705 79.795 57.715 ;
        RECT 84.760 57.705 85.130 57.715 ;
        RECT 90.085 57.705 90.455 57.715 ;
        RECT 95.420 57.705 95.790 57.715 ;
        RECT 100.745 57.705 101.115 57.715 ;
        RECT 106.080 57.705 106.450 57.715 ;
        RECT 111.405 57.705 111.775 57.715 ;
        RECT 116.740 57.705 117.110 57.715 ;
        RECT 28.035 56.395 28.315 56.765 ;
        RECT 28.085 53.145 28.265 56.395 ;
        RECT 28.035 52.775 28.315 53.145 ;
        RECT 28.085 50.525 28.265 52.775 ;
        RECT 28.465 51.855 28.645 57.690 ;
        RECT 36.785 57.445 37.810 57.705 ;
        RECT 41.285 57.610 41.655 57.620 ;
        RECT 36.785 57.435 37.155 57.445 ;
        RECT 40.630 57.350 41.655 57.610 ;
        RECT 42.120 57.445 43.145 57.705 ;
        RECT 46.620 57.610 46.990 57.620 ;
        RECT 42.120 57.435 42.490 57.445 ;
        RECT 45.965 57.350 46.990 57.610 ;
        RECT 47.445 57.445 48.470 57.705 ;
        RECT 51.945 57.610 52.315 57.620 ;
        RECT 47.445 57.435 47.815 57.445 ;
        RECT 51.290 57.350 52.315 57.610 ;
        RECT 52.780 57.445 53.805 57.705 ;
        RECT 57.280 57.610 57.650 57.620 ;
        RECT 52.780 57.435 53.150 57.445 ;
        RECT 56.625 57.350 57.650 57.610 ;
        RECT 58.105 57.445 59.130 57.705 ;
        RECT 62.605 57.610 62.975 57.620 ;
        RECT 58.105 57.435 58.475 57.445 ;
        RECT 61.950 57.350 62.975 57.610 ;
        RECT 63.440 57.445 64.465 57.705 ;
        RECT 67.940 57.610 68.310 57.620 ;
        RECT 63.440 57.435 63.810 57.445 ;
        RECT 67.285 57.350 68.310 57.610 ;
        RECT 68.765 57.445 69.790 57.705 ;
        RECT 73.265 57.610 73.635 57.620 ;
        RECT 68.765 57.435 69.135 57.445 ;
        RECT 72.610 57.350 73.635 57.610 ;
        RECT 74.100 57.445 75.125 57.705 ;
        RECT 78.600 57.610 78.970 57.620 ;
        RECT 74.100 57.435 74.470 57.445 ;
        RECT 77.945 57.350 78.970 57.610 ;
        RECT 79.425 57.445 80.450 57.705 ;
        RECT 83.925 57.610 84.295 57.620 ;
        RECT 79.425 57.435 79.795 57.445 ;
        RECT 83.270 57.350 84.295 57.610 ;
        RECT 84.760 57.445 85.785 57.705 ;
        RECT 89.260 57.610 89.630 57.620 ;
        RECT 84.760 57.435 85.130 57.445 ;
        RECT 88.605 57.350 89.630 57.610 ;
        RECT 90.085 57.445 91.110 57.705 ;
        RECT 94.585 57.610 94.955 57.620 ;
        RECT 90.085 57.435 90.455 57.445 ;
        RECT 93.930 57.350 94.955 57.610 ;
        RECT 95.420 57.445 96.445 57.705 ;
        RECT 99.920 57.610 100.290 57.620 ;
        RECT 95.420 57.435 95.790 57.445 ;
        RECT 99.265 57.350 100.290 57.610 ;
        RECT 100.745 57.445 101.770 57.705 ;
        RECT 105.245 57.610 105.615 57.620 ;
        RECT 100.745 57.435 101.115 57.445 ;
        RECT 104.590 57.350 105.615 57.610 ;
        RECT 106.080 57.445 107.105 57.705 ;
        RECT 110.580 57.610 110.950 57.620 ;
        RECT 106.080 57.435 106.450 57.445 ;
        RECT 109.925 57.350 110.950 57.610 ;
        RECT 111.405 57.445 112.430 57.705 ;
        RECT 115.905 57.610 116.275 57.620 ;
        RECT 111.405 57.435 111.775 57.445 ;
        RECT 115.250 57.350 116.275 57.610 ;
        RECT 116.740 57.445 117.765 57.705 ;
        RECT 121.240 57.610 121.610 57.620 ;
        RECT 116.740 57.435 117.110 57.445 ;
        RECT 120.585 57.350 121.610 57.610 ;
        RECT 41.285 57.340 41.655 57.350 ;
        RECT 46.620 57.340 46.990 57.350 ;
        RECT 51.945 57.340 52.315 57.350 ;
        RECT 57.280 57.340 57.650 57.350 ;
        RECT 62.605 57.340 62.975 57.350 ;
        RECT 67.940 57.340 68.310 57.350 ;
        RECT 73.265 57.340 73.635 57.350 ;
        RECT 78.600 57.340 78.970 57.350 ;
        RECT 83.925 57.340 84.295 57.350 ;
        RECT 89.260 57.340 89.630 57.350 ;
        RECT 94.585 57.340 94.955 57.350 ;
        RECT 99.920 57.340 100.290 57.350 ;
        RECT 105.245 57.340 105.615 57.350 ;
        RECT 110.580 57.340 110.950 57.350 ;
        RECT 115.905 57.340 116.275 57.350 ;
        RECT 121.240 57.340 121.610 57.350 ;
        RECT 34.005 57.055 34.400 57.060 ;
        RECT 33.390 56.775 35.160 57.055 ;
        RECT 38.715 56.775 39.110 57.055 ;
        RECT 39.330 56.780 39.725 57.060 ;
        RECT 39.385 56.550 39.645 56.780 ;
        RECT 40.030 56.775 40.485 57.055 ;
        RECT 44.050 56.775 44.445 57.055 ;
        RECT 44.665 56.780 45.060 57.060 ;
        RECT 44.720 56.550 44.980 56.780 ;
        RECT 45.365 56.775 45.820 57.055 ;
        RECT 49.375 56.775 49.770 57.055 ;
        RECT 49.990 56.780 50.385 57.060 ;
        RECT 50.045 56.550 50.305 56.780 ;
        RECT 50.690 56.775 51.145 57.055 ;
        RECT 54.710 56.775 55.105 57.055 ;
        RECT 55.325 56.780 55.720 57.060 ;
        RECT 55.380 56.550 55.640 56.780 ;
        RECT 56.025 56.775 56.480 57.055 ;
        RECT 60.035 56.775 60.430 57.055 ;
        RECT 60.650 56.780 61.045 57.060 ;
        RECT 60.705 56.550 60.965 56.780 ;
        RECT 61.350 56.775 61.805 57.055 ;
        RECT 65.370 56.775 65.765 57.055 ;
        RECT 65.985 56.780 66.380 57.060 ;
        RECT 66.040 56.550 66.300 56.780 ;
        RECT 66.685 56.775 67.140 57.055 ;
        RECT 70.695 56.775 71.090 57.055 ;
        RECT 71.310 56.780 71.705 57.060 ;
        RECT 71.365 56.550 71.625 56.780 ;
        RECT 72.010 56.775 72.465 57.055 ;
        RECT 76.030 56.775 76.425 57.055 ;
        RECT 76.645 56.780 77.040 57.060 ;
        RECT 76.700 56.550 76.960 56.780 ;
        RECT 77.345 56.775 77.800 57.055 ;
        RECT 81.355 56.775 81.750 57.055 ;
        RECT 81.970 56.780 82.365 57.060 ;
        RECT 82.025 56.550 82.285 56.780 ;
        RECT 82.670 56.775 83.125 57.055 ;
        RECT 86.690 56.775 87.085 57.055 ;
        RECT 87.305 56.780 87.700 57.060 ;
        RECT 87.360 56.550 87.620 56.780 ;
        RECT 88.005 56.775 88.460 57.055 ;
        RECT 92.015 56.775 92.410 57.055 ;
        RECT 92.630 56.780 93.025 57.060 ;
        RECT 92.685 56.550 92.945 56.780 ;
        RECT 93.330 56.775 93.785 57.055 ;
        RECT 97.350 56.775 97.745 57.055 ;
        RECT 97.965 56.780 98.360 57.060 ;
        RECT 98.020 56.550 98.280 56.780 ;
        RECT 98.665 56.775 99.120 57.055 ;
        RECT 102.675 56.775 103.070 57.055 ;
        RECT 103.290 56.780 103.685 57.060 ;
        RECT 103.345 56.550 103.605 56.780 ;
        RECT 103.990 56.775 104.445 57.055 ;
        RECT 108.010 56.775 108.405 57.055 ;
        RECT 108.625 56.780 109.020 57.060 ;
        RECT 108.680 56.550 108.940 56.780 ;
        RECT 109.325 56.775 109.780 57.055 ;
        RECT 113.335 56.775 113.730 57.055 ;
        RECT 113.950 56.780 114.345 57.060 ;
        RECT 114.005 56.550 114.265 56.780 ;
        RECT 114.650 56.775 115.105 57.055 ;
        RECT 118.670 56.775 119.065 57.055 ;
        RECT 119.285 56.780 119.680 57.060 ;
        RECT 124.610 57.055 125.005 57.060 ;
        RECT 119.340 56.550 119.600 56.780 ;
        RECT 119.985 56.775 120.440 57.055 ;
        RECT 123.995 56.775 125.765 57.055 ;
        RECT 36.785 56.405 37.155 56.415 ;
        RECT 36.785 56.145 37.860 56.405 ;
        RECT 39.385 56.270 41.015 56.550 ;
        RECT 42.120 56.405 42.490 56.415 ;
        RECT 42.120 56.145 43.195 56.405 ;
        RECT 44.720 56.270 46.350 56.550 ;
        RECT 47.445 56.405 47.815 56.415 ;
        RECT 47.445 56.145 48.520 56.405 ;
        RECT 50.045 56.270 51.675 56.550 ;
        RECT 52.780 56.405 53.150 56.415 ;
        RECT 52.780 56.145 53.855 56.405 ;
        RECT 55.380 56.270 57.010 56.550 ;
        RECT 58.105 56.405 58.475 56.415 ;
        RECT 58.105 56.145 59.180 56.405 ;
        RECT 60.705 56.270 62.335 56.550 ;
        RECT 63.440 56.405 63.810 56.415 ;
        RECT 63.440 56.145 64.515 56.405 ;
        RECT 66.040 56.270 67.670 56.550 ;
        RECT 68.765 56.405 69.135 56.415 ;
        RECT 68.765 56.145 69.840 56.405 ;
        RECT 71.365 56.270 72.995 56.550 ;
        RECT 74.100 56.405 74.470 56.415 ;
        RECT 74.100 56.145 75.175 56.405 ;
        RECT 76.700 56.270 78.330 56.550 ;
        RECT 79.425 56.405 79.795 56.415 ;
        RECT 79.425 56.145 80.500 56.405 ;
        RECT 82.025 56.270 83.655 56.550 ;
        RECT 84.760 56.405 85.130 56.415 ;
        RECT 84.760 56.145 85.835 56.405 ;
        RECT 87.360 56.270 88.990 56.550 ;
        RECT 90.085 56.405 90.455 56.415 ;
        RECT 90.085 56.145 91.160 56.405 ;
        RECT 92.685 56.270 94.315 56.550 ;
        RECT 95.420 56.405 95.790 56.415 ;
        RECT 95.420 56.145 96.495 56.405 ;
        RECT 98.020 56.270 99.650 56.550 ;
        RECT 100.745 56.405 101.115 56.415 ;
        RECT 100.745 56.145 101.820 56.405 ;
        RECT 103.345 56.270 104.975 56.550 ;
        RECT 106.080 56.405 106.450 56.415 ;
        RECT 106.080 56.145 107.155 56.405 ;
        RECT 108.680 56.270 110.310 56.550 ;
        RECT 111.405 56.405 111.775 56.415 ;
        RECT 111.405 56.145 112.480 56.405 ;
        RECT 114.005 56.270 115.635 56.550 ;
        RECT 116.740 56.405 117.110 56.415 ;
        RECT 116.740 56.145 117.815 56.405 ;
        RECT 119.340 56.270 120.970 56.550 ;
        RECT 36.785 56.135 37.155 56.145 ;
        RECT 42.120 56.135 42.490 56.145 ;
        RECT 47.445 56.135 47.815 56.145 ;
        RECT 52.780 56.135 53.150 56.145 ;
        RECT 58.105 56.135 58.475 56.145 ;
        RECT 63.440 56.135 63.810 56.145 ;
        RECT 68.765 56.135 69.135 56.145 ;
        RECT 74.100 56.135 74.470 56.145 ;
        RECT 79.425 56.135 79.795 56.145 ;
        RECT 84.760 56.135 85.130 56.145 ;
        RECT 90.085 56.135 90.455 56.145 ;
        RECT 95.420 56.135 95.790 56.145 ;
        RECT 100.745 56.135 101.115 56.145 ;
        RECT 106.080 56.135 106.450 56.145 ;
        RECT 111.405 56.135 111.775 56.145 ;
        RECT 116.740 56.135 117.110 56.145 ;
        RECT 41.290 55.775 41.660 55.785 ;
        RECT 46.625 55.775 46.995 55.785 ;
        RECT 51.950 55.775 52.320 55.785 ;
        RECT 57.285 55.775 57.655 55.785 ;
        RECT 62.610 55.775 62.980 55.785 ;
        RECT 67.945 55.775 68.315 55.785 ;
        RECT 73.270 55.775 73.640 55.785 ;
        RECT 78.605 55.775 78.975 55.785 ;
        RECT 83.930 55.775 84.300 55.785 ;
        RECT 89.265 55.775 89.635 55.785 ;
        RECT 94.590 55.775 94.960 55.785 ;
        RECT 99.925 55.775 100.295 55.785 ;
        RECT 105.250 55.775 105.620 55.785 ;
        RECT 110.585 55.775 110.955 55.785 ;
        RECT 115.910 55.775 116.280 55.785 ;
        RECT 121.245 55.775 121.615 55.785 ;
        RECT 40.630 55.515 41.660 55.775 ;
        RECT 45.965 55.515 46.995 55.775 ;
        RECT 51.290 55.515 52.320 55.775 ;
        RECT 56.625 55.515 57.655 55.775 ;
        RECT 61.950 55.515 62.980 55.775 ;
        RECT 67.285 55.515 68.315 55.775 ;
        RECT 72.610 55.515 73.640 55.775 ;
        RECT 77.945 55.515 78.975 55.775 ;
        RECT 83.270 55.515 84.300 55.775 ;
        RECT 88.605 55.515 89.635 55.775 ;
        RECT 93.930 55.515 94.960 55.775 ;
        RECT 99.265 55.515 100.295 55.775 ;
        RECT 104.590 55.515 105.620 55.775 ;
        RECT 109.925 55.515 110.955 55.775 ;
        RECT 115.250 55.515 116.280 55.775 ;
        RECT 120.585 55.515 121.615 55.775 ;
        RECT 41.290 55.505 41.660 55.515 ;
        RECT 46.625 55.505 46.995 55.515 ;
        RECT 51.950 55.505 52.320 55.515 ;
        RECT 57.285 55.505 57.655 55.515 ;
        RECT 62.610 55.505 62.980 55.515 ;
        RECT 67.945 55.505 68.315 55.515 ;
        RECT 73.270 55.505 73.640 55.515 ;
        RECT 78.605 55.505 78.975 55.515 ;
        RECT 83.930 55.505 84.300 55.515 ;
        RECT 89.265 55.505 89.635 55.515 ;
        RECT 94.590 55.505 94.960 55.515 ;
        RECT 99.925 55.505 100.295 55.515 ;
        RECT 105.250 55.505 105.620 55.515 ;
        RECT 110.585 55.505 110.955 55.515 ;
        RECT 115.910 55.505 116.280 55.515 ;
        RECT 121.245 55.505 121.615 55.515 ;
        RECT 36.790 54.040 37.160 54.050 ;
        RECT 42.125 54.040 42.495 54.050 ;
        RECT 47.450 54.040 47.820 54.050 ;
        RECT 52.785 54.040 53.155 54.050 ;
        RECT 58.110 54.040 58.480 54.050 ;
        RECT 63.445 54.040 63.815 54.050 ;
        RECT 68.770 54.040 69.140 54.050 ;
        RECT 74.105 54.040 74.475 54.050 ;
        RECT 79.430 54.040 79.800 54.050 ;
        RECT 84.765 54.040 85.135 54.050 ;
        RECT 90.090 54.040 90.460 54.050 ;
        RECT 95.425 54.040 95.795 54.050 ;
        RECT 100.750 54.040 101.120 54.050 ;
        RECT 106.085 54.040 106.455 54.050 ;
        RECT 111.410 54.040 111.780 54.050 ;
        RECT 116.745 54.040 117.115 54.050 ;
        RECT 36.790 53.780 37.810 54.040 ;
        RECT 42.125 53.780 43.145 54.040 ;
        RECT 47.450 53.780 48.470 54.040 ;
        RECT 52.785 53.780 53.805 54.040 ;
        RECT 58.110 53.780 59.130 54.040 ;
        RECT 63.445 53.780 64.465 54.040 ;
        RECT 68.770 53.780 69.790 54.040 ;
        RECT 74.105 53.780 75.125 54.040 ;
        RECT 79.430 53.780 80.450 54.040 ;
        RECT 84.765 53.780 85.785 54.040 ;
        RECT 90.090 53.780 91.110 54.040 ;
        RECT 95.425 53.780 96.445 54.040 ;
        RECT 100.750 53.780 101.770 54.040 ;
        RECT 106.085 53.780 107.105 54.040 ;
        RECT 111.410 53.780 112.430 54.040 ;
        RECT 116.745 53.780 117.765 54.040 ;
        RECT 36.790 53.770 37.160 53.780 ;
        RECT 42.125 53.770 42.495 53.780 ;
        RECT 47.450 53.770 47.820 53.780 ;
        RECT 52.785 53.770 53.155 53.780 ;
        RECT 58.110 53.770 58.480 53.780 ;
        RECT 63.445 53.770 63.815 53.780 ;
        RECT 68.770 53.770 69.140 53.780 ;
        RECT 74.105 53.770 74.475 53.780 ;
        RECT 79.430 53.770 79.800 53.780 ;
        RECT 84.765 53.770 85.135 53.780 ;
        RECT 90.090 53.770 90.460 53.780 ;
        RECT 95.425 53.770 95.795 53.780 ;
        RECT 100.750 53.770 101.120 53.780 ;
        RECT 106.085 53.770 106.455 53.780 ;
        RECT 111.410 53.770 111.780 53.780 ;
        RECT 116.745 53.770 117.115 53.780 ;
        RECT 41.285 53.390 41.655 53.400 ;
        RECT 46.620 53.390 46.990 53.400 ;
        RECT 51.945 53.390 52.315 53.400 ;
        RECT 57.280 53.390 57.650 53.400 ;
        RECT 62.605 53.390 62.975 53.400 ;
        RECT 67.940 53.390 68.310 53.400 ;
        RECT 73.265 53.390 73.635 53.400 ;
        RECT 78.600 53.390 78.970 53.400 ;
        RECT 83.925 53.390 84.295 53.400 ;
        RECT 89.260 53.390 89.630 53.400 ;
        RECT 94.585 53.390 94.955 53.400 ;
        RECT 99.920 53.390 100.290 53.400 ;
        RECT 105.245 53.390 105.615 53.400 ;
        RECT 110.580 53.390 110.950 53.400 ;
        RECT 115.905 53.390 116.275 53.400 ;
        RECT 121.240 53.390 121.610 53.400 ;
        RECT 37.430 52.995 39.055 53.275 ;
        RECT 40.580 53.130 41.655 53.390 ;
        RECT 41.285 53.120 41.655 53.130 ;
        RECT 42.765 52.995 44.390 53.275 ;
        RECT 45.915 53.130 46.990 53.390 ;
        RECT 46.620 53.120 46.990 53.130 ;
        RECT 48.090 52.995 49.715 53.275 ;
        RECT 51.240 53.130 52.315 53.390 ;
        RECT 51.945 53.120 52.315 53.130 ;
        RECT 53.425 52.995 55.050 53.275 ;
        RECT 56.575 53.130 57.650 53.390 ;
        RECT 57.280 53.120 57.650 53.130 ;
        RECT 58.750 52.995 60.375 53.275 ;
        RECT 61.900 53.130 62.975 53.390 ;
        RECT 62.605 53.120 62.975 53.130 ;
        RECT 64.085 52.995 65.710 53.275 ;
        RECT 67.235 53.130 68.310 53.390 ;
        RECT 67.940 53.120 68.310 53.130 ;
        RECT 69.410 52.995 71.035 53.275 ;
        RECT 72.560 53.130 73.635 53.390 ;
        RECT 73.265 53.120 73.635 53.130 ;
        RECT 74.745 52.995 76.370 53.275 ;
        RECT 77.895 53.130 78.970 53.390 ;
        RECT 78.600 53.120 78.970 53.130 ;
        RECT 80.070 52.995 81.695 53.275 ;
        RECT 83.220 53.130 84.295 53.390 ;
        RECT 83.925 53.120 84.295 53.130 ;
        RECT 85.405 52.995 87.030 53.275 ;
        RECT 88.555 53.130 89.630 53.390 ;
        RECT 89.260 53.120 89.630 53.130 ;
        RECT 90.730 52.995 92.355 53.275 ;
        RECT 93.880 53.130 94.955 53.390 ;
        RECT 94.585 53.120 94.955 53.130 ;
        RECT 96.065 52.995 97.690 53.275 ;
        RECT 99.215 53.130 100.290 53.390 ;
        RECT 99.920 53.120 100.290 53.130 ;
        RECT 101.390 52.995 103.015 53.275 ;
        RECT 104.540 53.130 105.615 53.390 ;
        RECT 105.245 53.120 105.615 53.130 ;
        RECT 106.725 52.995 108.350 53.275 ;
        RECT 109.875 53.130 110.950 53.390 ;
        RECT 110.580 53.120 110.950 53.130 ;
        RECT 112.050 52.995 113.675 53.275 ;
        RECT 115.200 53.130 116.275 53.390 ;
        RECT 115.905 53.120 116.275 53.130 ;
        RECT 117.385 52.995 119.010 53.275 ;
        RECT 120.535 53.130 121.610 53.390 ;
        RECT 121.240 53.120 121.610 53.130 ;
        RECT 38.795 52.695 39.055 52.995 ;
        RECT 44.130 52.695 44.390 52.995 ;
        RECT 49.455 52.695 49.715 52.995 ;
        RECT 54.790 52.695 55.050 52.995 ;
        RECT 60.115 52.695 60.375 52.995 ;
        RECT 65.450 52.695 65.710 52.995 ;
        RECT 70.775 52.695 71.035 52.995 ;
        RECT 76.110 52.695 76.370 52.995 ;
        RECT 81.435 52.695 81.695 52.995 ;
        RECT 86.770 52.695 87.030 52.995 ;
        RECT 92.095 52.695 92.355 52.995 ;
        RECT 97.430 52.695 97.690 52.995 ;
        RECT 102.755 52.695 103.015 52.995 ;
        RECT 108.090 52.695 108.350 52.995 ;
        RECT 113.415 52.695 113.675 52.995 ;
        RECT 118.750 52.695 119.010 52.995 ;
        RECT 32.625 52.415 34.390 52.695 ;
        RECT 37.950 52.415 38.485 52.695 ;
        RECT 38.715 52.415 39.110 52.695 ;
        RECT 39.330 52.415 39.730 52.695 ;
        RECT 43.285 52.415 43.820 52.695 ;
        RECT 44.050 52.415 44.445 52.695 ;
        RECT 44.665 52.415 45.065 52.695 ;
        RECT 48.610 52.415 49.145 52.695 ;
        RECT 49.375 52.415 49.770 52.695 ;
        RECT 49.990 52.415 50.390 52.695 ;
        RECT 53.945 52.415 54.480 52.695 ;
        RECT 54.710 52.415 55.105 52.695 ;
        RECT 55.325 52.415 55.725 52.695 ;
        RECT 59.270 52.415 59.805 52.695 ;
        RECT 60.035 52.415 60.430 52.695 ;
        RECT 60.650 52.415 61.050 52.695 ;
        RECT 64.605 52.415 65.140 52.695 ;
        RECT 65.370 52.415 65.765 52.695 ;
        RECT 65.985 52.415 66.385 52.695 ;
        RECT 69.930 52.415 70.465 52.695 ;
        RECT 70.695 52.415 71.090 52.695 ;
        RECT 71.310 52.415 71.710 52.695 ;
        RECT 75.265 52.415 75.800 52.695 ;
        RECT 76.030 52.415 76.425 52.695 ;
        RECT 76.645 52.415 77.045 52.695 ;
        RECT 80.590 52.415 81.125 52.695 ;
        RECT 81.355 52.415 81.750 52.695 ;
        RECT 81.970 52.415 82.370 52.695 ;
        RECT 85.925 52.415 86.460 52.695 ;
        RECT 86.690 52.415 87.085 52.695 ;
        RECT 87.305 52.415 87.705 52.695 ;
        RECT 91.250 52.415 91.785 52.695 ;
        RECT 92.015 52.415 92.410 52.695 ;
        RECT 92.630 52.415 93.030 52.695 ;
        RECT 96.585 52.415 97.120 52.695 ;
        RECT 97.350 52.415 97.745 52.695 ;
        RECT 97.965 52.415 98.365 52.695 ;
        RECT 101.910 52.415 102.445 52.695 ;
        RECT 102.675 52.415 103.070 52.695 ;
        RECT 103.290 52.415 103.690 52.695 ;
        RECT 107.245 52.415 107.780 52.695 ;
        RECT 108.010 52.415 108.405 52.695 ;
        RECT 108.625 52.415 109.025 52.695 ;
        RECT 112.570 52.415 113.105 52.695 ;
        RECT 113.335 52.415 113.730 52.695 ;
        RECT 113.950 52.415 114.350 52.695 ;
        RECT 117.905 52.415 118.440 52.695 ;
        RECT 118.670 52.415 119.065 52.695 ;
        RECT 119.285 52.415 119.685 52.695 ;
        RECT 123.230 52.415 124.995 52.695 ;
        RECT 36.785 52.195 37.155 52.205 ;
        RECT 42.120 52.195 42.490 52.205 ;
        RECT 47.445 52.195 47.815 52.205 ;
        RECT 52.780 52.195 53.150 52.205 ;
        RECT 58.105 52.195 58.475 52.205 ;
        RECT 63.440 52.195 63.810 52.205 ;
        RECT 68.765 52.195 69.135 52.205 ;
        RECT 74.100 52.195 74.470 52.205 ;
        RECT 79.425 52.195 79.795 52.205 ;
        RECT 84.760 52.195 85.130 52.205 ;
        RECT 90.085 52.195 90.455 52.205 ;
        RECT 95.420 52.195 95.790 52.205 ;
        RECT 100.745 52.195 101.115 52.205 ;
        RECT 106.080 52.195 106.450 52.205 ;
        RECT 111.405 52.195 111.775 52.205 ;
        RECT 116.740 52.195 117.110 52.205 ;
        RECT 36.785 51.935 37.810 52.195 ;
        RECT 41.285 52.105 41.655 52.115 ;
        RECT 36.785 51.925 37.155 51.935 ;
        RECT 28.415 51.485 28.695 51.855 ;
        RECT 40.630 51.845 41.655 52.105 ;
        RECT 42.120 51.935 43.145 52.195 ;
        RECT 46.620 52.105 46.990 52.115 ;
        RECT 42.120 51.925 42.490 51.935 ;
        RECT 45.965 51.845 46.990 52.105 ;
        RECT 47.445 51.935 48.470 52.195 ;
        RECT 51.945 52.105 52.315 52.115 ;
        RECT 47.445 51.925 47.815 51.935 ;
        RECT 51.290 51.845 52.315 52.105 ;
        RECT 52.780 51.935 53.805 52.195 ;
        RECT 57.280 52.105 57.650 52.115 ;
        RECT 52.780 51.925 53.150 51.935 ;
        RECT 56.625 51.845 57.650 52.105 ;
        RECT 58.105 51.935 59.130 52.195 ;
        RECT 62.605 52.105 62.975 52.115 ;
        RECT 58.105 51.925 58.475 51.935 ;
        RECT 61.950 51.845 62.975 52.105 ;
        RECT 63.440 51.935 64.465 52.195 ;
        RECT 67.940 52.105 68.310 52.115 ;
        RECT 63.440 51.925 63.810 51.935 ;
        RECT 67.285 51.845 68.310 52.105 ;
        RECT 68.765 51.935 69.790 52.195 ;
        RECT 73.265 52.105 73.635 52.115 ;
        RECT 68.765 51.925 69.135 51.935 ;
        RECT 72.610 51.845 73.635 52.105 ;
        RECT 74.100 51.935 75.125 52.195 ;
        RECT 78.600 52.105 78.970 52.115 ;
        RECT 74.100 51.925 74.470 51.935 ;
        RECT 77.945 51.845 78.970 52.105 ;
        RECT 79.425 51.935 80.450 52.195 ;
        RECT 83.925 52.105 84.295 52.115 ;
        RECT 79.425 51.925 79.795 51.935 ;
        RECT 83.270 51.845 84.295 52.105 ;
        RECT 84.760 51.935 85.785 52.195 ;
        RECT 89.260 52.105 89.630 52.115 ;
        RECT 84.760 51.925 85.130 51.935 ;
        RECT 88.605 51.845 89.630 52.105 ;
        RECT 90.085 51.935 91.110 52.195 ;
        RECT 94.585 52.105 94.955 52.115 ;
        RECT 90.085 51.925 90.455 51.935 ;
        RECT 93.930 51.845 94.955 52.105 ;
        RECT 95.420 51.935 96.445 52.195 ;
        RECT 99.920 52.105 100.290 52.115 ;
        RECT 95.420 51.925 95.790 51.935 ;
        RECT 99.265 51.845 100.290 52.105 ;
        RECT 100.745 51.935 101.770 52.195 ;
        RECT 105.245 52.105 105.615 52.115 ;
        RECT 100.745 51.925 101.115 51.935 ;
        RECT 104.590 51.845 105.615 52.105 ;
        RECT 106.080 51.935 107.105 52.195 ;
        RECT 110.580 52.105 110.950 52.115 ;
        RECT 106.080 51.925 106.450 51.935 ;
        RECT 109.925 51.845 110.950 52.105 ;
        RECT 111.405 51.935 112.430 52.195 ;
        RECT 115.905 52.105 116.275 52.115 ;
        RECT 111.405 51.925 111.775 51.935 ;
        RECT 115.250 51.845 116.275 52.105 ;
        RECT 116.740 51.935 117.765 52.195 ;
        RECT 121.240 52.105 121.610 52.115 ;
        RECT 116.740 51.925 117.110 51.935 ;
        RECT 120.585 51.845 121.610 52.105 ;
        RECT 41.285 51.835 41.655 51.845 ;
        RECT 46.620 51.835 46.990 51.845 ;
        RECT 51.945 51.835 52.315 51.845 ;
        RECT 57.280 51.835 57.650 51.845 ;
        RECT 62.605 51.835 62.975 51.845 ;
        RECT 67.940 51.835 68.310 51.845 ;
        RECT 73.265 51.835 73.635 51.845 ;
        RECT 78.600 51.835 78.970 51.845 ;
        RECT 83.925 51.835 84.295 51.845 ;
        RECT 89.260 51.835 89.630 51.845 ;
        RECT 94.585 51.835 94.955 51.845 ;
        RECT 99.920 51.835 100.290 51.845 ;
        RECT 105.245 51.835 105.615 51.845 ;
        RECT 110.580 51.835 110.950 51.845 ;
        RECT 115.905 51.835 116.275 51.845 ;
        RECT 121.240 51.835 121.610 51.845 ;
        RECT 28.030 50.155 28.310 50.525 ;
        RECT 27.655 49.505 27.935 49.875 ;
        RECT 27.275 48.215 27.555 48.585 ;
        RECT 27.325 44.965 27.505 48.215 ;
        RECT 27.705 46.255 27.885 49.505 ;
        RECT 27.650 45.885 27.930 46.255 ;
        RECT 27.275 44.595 27.555 44.965 ;
        RECT 27.325 34.805 27.505 44.595 ;
        RECT 27.275 34.435 27.555 34.805 ;
        RECT 27.325 31.185 27.505 34.435 ;
        RECT 27.705 33.515 27.885 45.885 ;
        RECT 28.085 44.320 28.265 50.155 ;
        RECT 28.465 49.230 28.645 51.485 ;
        RECT 36.785 50.170 37.155 50.180 ;
        RECT 42.120 50.170 42.490 50.180 ;
        RECT 47.445 50.170 47.815 50.180 ;
        RECT 52.780 50.170 53.150 50.180 ;
        RECT 58.105 50.170 58.475 50.180 ;
        RECT 63.440 50.170 63.810 50.180 ;
        RECT 68.765 50.170 69.135 50.180 ;
        RECT 74.100 50.170 74.470 50.180 ;
        RECT 79.425 50.170 79.795 50.180 ;
        RECT 84.760 50.170 85.130 50.180 ;
        RECT 90.085 50.170 90.455 50.180 ;
        RECT 95.420 50.170 95.790 50.180 ;
        RECT 100.745 50.170 101.115 50.180 ;
        RECT 106.080 50.170 106.450 50.180 ;
        RECT 111.405 50.170 111.775 50.180 ;
        RECT 116.740 50.170 117.110 50.180 ;
        RECT 36.785 49.910 37.810 50.170 ;
        RECT 41.285 50.075 41.655 50.085 ;
        RECT 36.785 49.900 37.155 49.910 ;
        RECT 40.630 49.815 41.655 50.075 ;
        RECT 42.120 49.910 43.145 50.170 ;
        RECT 46.620 50.075 46.990 50.085 ;
        RECT 42.120 49.900 42.490 49.910 ;
        RECT 45.965 49.815 46.990 50.075 ;
        RECT 47.445 49.910 48.470 50.170 ;
        RECT 51.945 50.075 52.315 50.085 ;
        RECT 47.445 49.900 47.815 49.910 ;
        RECT 51.290 49.815 52.315 50.075 ;
        RECT 52.780 49.910 53.805 50.170 ;
        RECT 57.280 50.075 57.650 50.085 ;
        RECT 52.780 49.900 53.150 49.910 ;
        RECT 56.625 49.815 57.650 50.075 ;
        RECT 58.105 49.910 59.130 50.170 ;
        RECT 62.605 50.075 62.975 50.085 ;
        RECT 58.105 49.900 58.475 49.910 ;
        RECT 61.950 49.815 62.975 50.075 ;
        RECT 63.440 49.910 64.465 50.170 ;
        RECT 67.940 50.075 68.310 50.085 ;
        RECT 63.440 49.900 63.810 49.910 ;
        RECT 67.285 49.815 68.310 50.075 ;
        RECT 68.765 49.910 69.790 50.170 ;
        RECT 73.265 50.075 73.635 50.085 ;
        RECT 68.765 49.900 69.135 49.910 ;
        RECT 72.610 49.815 73.635 50.075 ;
        RECT 74.100 49.910 75.125 50.170 ;
        RECT 78.600 50.075 78.970 50.085 ;
        RECT 74.100 49.900 74.470 49.910 ;
        RECT 77.945 49.815 78.970 50.075 ;
        RECT 79.425 49.910 80.450 50.170 ;
        RECT 83.925 50.075 84.295 50.085 ;
        RECT 79.425 49.900 79.795 49.910 ;
        RECT 83.270 49.815 84.295 50.075 ;
        RECT 84.760 49.910 85.785 50.170 ;
        RECT 89.260 50.075 89.630 50.085 ;
        RECT 84.760 49.900 85.130 49.910 ;
        RECT 88.605 49.815 89.630 50.075 ;
        RECT 90.085 49.910 91.110 50.170 ;
        RECT 94.585 50.075 94.955 50.085 ;
        RECT 90.085 49.900 90.455 49.910 ;
        RECT 93.930 49.815 94.955 50.075 ;
        RECT 95.420 49.910 96.445 50.170 ;
        RECT 99.920 50.075 100.290 50.085 ;
        RECT 95.420 49.900 95.790 49.910 ;
        RECT 99.265 49.815 100.290 50.075 ;
        RECT 100.745 49.910 101.770 50.170 ;
        RECT 105.245 50.075 105.615 50.085 ;
        RECT 100.745 49.900 101.115 49.910 ;
        RECT 104.590 49.815 105.615 50.075 ;
        RECT 106.080 49.910 107.105 50.170 ;
        RECT 110.580 50.075 110.950 50.085 ;
        RECT 106.080 49.900 106.450 49.910 ;
        RECT 109.925 49.815 110.950 50.075 ;
        RECT 111.405 49.910 112.430 50.170 ;
        RECT 115.905 50.075 116.275 50.085 ;
        RECT 111.405 49.900 111.775 49.910 ;
        RECT 115.250 49.815 116.275 50.075 ;
        RECT 116.740 49.910 117.765 50.170 ;
        RECT 121.240 50.075 121.610 50.085 ;
        RECT 116.740 49.900 117.110 49.910 ;
        RECT 120.585 49.815 121.610 50.075 ;
        RECT 41.285 49.805 41.655 49.815 ;
        RECT 46.620 49.805 46.990 49.815 ;
        RECT 51.945 49.805 52.315 49.815 ;
        RECT 57.280 49.805 57.650 49.815 ;
        RECT 62.605 49.805 62.975 49.815 ;
        RECT 67.940 49.805 68.310 49.815 ;
        RECT 73.265 49.805 73.635 49.815 ;
        RECT 78.600 49.805 78.970 49.815 ;
        RECT 83.925 49.805 84.295 49.815 ;
        RECT 89.260 49.805 89.630 49.815 ;
        RECT 94.585 49.805 94.955 49.815 ;
        RECT 99.920 49.805 100.290 49.815 ;
        RECT 105.245 49.805 105.615 49.815 ;
        RECT 110.580 49.805 110.950 49.815 ;
        RECT 115.905 49.805 116.275 49.815 ;
        RECT 121.240 49.805 121.610 49.815 ;
        RECT 34.005 49.520 34.400 49.525 ;
        RECT 33.390 49.240 35.160 49.520 ;
        RECT 38.715 49.240 39.110 49.520 ;
        RECT 39.330 49.245 39.730 49.525 ;
        RECT 40.015 49.240 40.485 49.520 ;
        RECT 44.050 49.240 44.445 49.520 ;
        RECT 44.665 49.245 45.065 49.525 ;
        RECT 45.350 49.240 45.820 49.520 ;
        RECT 49.375 49.240 49.770 49.520 ;
        RECT 49.990 49.245 50.390 49.525 ;
        RECT 50.675 49.240 51.145 49.520 ;
        RECT 54.710 49.240 55.105 49.520 ;
        RECT 55.325 49.245 55.725 49.525 ;
        RECT 56.010 49.240 56.480 49.520 ;
        RECT 60.035 49.240 60.430 49.520 ;
        RECT 60.650 49.245 61.050 49.525 ;
        RECT 61.335 49.240 61.805 49.520 ;
        RECT 65.370 49.240 65.765 49.520 ;
        RECT 65.985 49.245 66.385 49.525 ;
        RECT 66.670 49.240 67.140 49.520 ;
        RECT 70.695 49.240 71.090 49.520 ;
        RECT 71.310 49.245 71.710 49.525 ;
        RECT 71.995 49.240 72.465 49.520 ;
        RECT 76.030 49.240 76.425 49.520 ;
        RECT 76.645 49.245 77.045 49.525 ;
        RECT 77.330 49.240 77.800 49.520 ;
        RECT 81.355 49.240 81.750 49.520 ;
        RECT 81.970 49.245 82.370 49.525 ;
        RECT 82.655 49.240 83.125 49.520 ;
        RECT 86.690 49.240 87.085 49.520 ;
        RECT 87.305 49.245 87.705 49.525 ;
        RECT 87.990 49.240 88.460 49.520 ;
        RECT 92.015 49.240 92.410 49.520 ;
        RECT 92.630 49.245 93.030 49.525 ;
        RECT 93.315 49.240 93.785 49.520 ;
        RECT 97.350 49.240 97.745 49.520 ;
        RECT 97.965 49.245 98.365 49.525 ;
        RECT 98.650 49.240 99.120 49.520 ;
        RECT 102.675 49.240 103.070 49.520 ;
        RECT 103.290 49.245 103.690 49.525 ;
        RECT 103.975 49.240 104.445 49.520 ;
        RECT 108.010 49.240 108.405 49.520 ;
        RECT 108.625 49.245 109.025 49.525 ;
        RECT 109.310 49.240 109.780 49.520 ;
        RECT 113.335 49.240 113.730 49.520 ;
        RECT 113.950 49.245 114.350 49.525 ;
        RECT 114.635 49.240 115.105 49.520 ;
        RECT 118.670 49.240 119.065 49.520 ;
        RECT 119.285 49.245 119.685 49.525 ;
        RECT 124.610 49.520 125.005 49.525 ;
        RECT 119.970 49.240 120.440 49.520 ;
        RECT 123.995 49.240 125.765 49.520 ;
        RECT 28.415 48.860 28.695 49.230 ;
        RECT 36.785 48.870 37.155 48.880 ;
        RECT 42.120 48.870 42.490 48.880 ;
        RECT 47.445 48.870 47.815 48.880 ;
        RECT 52.780 48.870 53.150 48.880 ;
        RECT 58.105 48.870 58.475 48.880 ;
        RECT 63.440 48.870 63.810 48.880 ;
        RECT 68.765 48.870 69.135 48.880 ;
        RECT 74.100 48.870 74.470 48.880 ;
        RECT 79.425 48.870 79.795 48.880 ;
        RECT 84.760 48.870 85.130 48.880 ;
        RECT 90.085 48.870 90.455 48.880 ;
        RECT 95.420 48.870 95.790 48.880 ;
        RECT 100.745 48.870 101.115 48.880 ;
        RECT 106.080 48.870 106.450 48.880 ;
        RECT 111.405 48.870 111.775 48.880 ;
        RECT 116.740 48.870 117.110 48.880 ;
        RECT 28.465 45.610 28.645 48.860 ;
        RECT 36.785 48.610 37.860 48.870 ;
        RECT 42.120 48.610 43.195 48.870 ;
        RECT 47.445 48.610 48.520 48.870 ;
        RECT 52.780 48.610 53.855 48.870 ;
        RECT 58.105 48.610 59.180 48.870 ;
        RECT 63.440 48.610 64.515 48.870 ;
        RECT 68.765 48.610 69.840 48.870 ;
        RECT 74.100 48.610 75.175 48.870 ;
        RECT 79.425 48.610 80.500 48.870 ;
        RECT 84.760 48.610 85.835 48.870 ;
        RECT 90.085 48.610 91.160 48.870 ;
        RECT 95.420 48.610 96.495 48.870 ;
        RECT 100.745 48.610 101.820 48.870 ;
        RECT 106.080 48.610 107.155 48.870 ;
        RECT 111.405 48.610 112.480 48.870 ;
        RECT 116.740 48.610 117.815 48.870 ;
        RECT 36.785 48.600 37.155 48.610 ;
        RECT 42.120 48.600 42.490 48.610 ;
        RECT 47.445 48.600 47.815 48.610 ;
        RECT 52.780 48.600 53.150 48.610 ;
        RECT 58.105 48.600 58.475 48.610 ;
        RECT 63.440 48.600 63.810 48.610 ;
        RECT 68.765 48.600 69.135 48.610 ;
        RECT 74.100 48.600 74.470 48.610 ;
        RECT 79.425 48.600 79.795 48.610 ;
        RECT 84.760 48.600 85.130 48.610 ;
        RECT 90.085 48.600 90.455 48.610 ;
        RECT 95.420 48.600 95.790 48.610 ;
        RECT 100.745 48.600 101.115 48.610 ;
        RECT 106.080 48.600 106.450 48.610 ;
        RECT 111.405 48.600 111.775 48.610 ;
        RECT 116.740 48.600 117.110 48.610 ;
        RECT 41.290 48.240 41.660 48.250 ;
        RECT 46.625 48.240 46.995 48.250 ;
        RECT 51.950 48.240 52.320 48.250 ;
        RECT 57.285 48.240 57.655 48.250 ;
        RECT 62.610 48.240 62.980 48.250 ;
        RECT 67.945 48.240 68.315 48.250 ;
        RECT 73.270 48.240 73.640 48.250 ;
        RECT 78.605 48.240 78.975 48.250 ;
        RECT 83.930 48.240 84.300 48.250 ;
        RECT 89.265 48.240 89.635 48.250 ;
        RECT 94.590 48.240 94.960 48.250 ;
        RECT 99.925 48.240 100.295 48.250 ;
        RECT 105.250 48.240 105.620 48.250 ;
        RECT 110.585 48.240 110.955 48.250 ;
        RECT 115.910 48.240 116.280 48.250 ;
        RECT 121.245 48.240 121.615 48.250 ;
        RECT 40.630 47.980 41.660 48.240 ;
        RECT 45.965 47.980 46.995 48.240 ;
        RECT 51.290 47.980 52.320 48.240 ;
        RECT 56.625 47.980 57.655 48.240 ;
        RECT 61.950 47.980 62.980 48.240 ;
        RECT 67.285 47.980 68.315 48.240 ;
        RECT 72.610 47.980 73.640 48.240 ;
        RECT 77.945 47.980 78.975 48.240 ;
        RECT 83.270 47.980 84.300 48.240 ;
        RECT 88.605 47.980 89.635 48.240 ;
        RECT 93.930 47.980 94.960 48.240 ;
        RECT 99.265 47.980 100.295 48.240 ;
        RECT 104.590 47.980 105.620 48.240 ;
        RECT 109.925 47.980 110.955 48.240 ;
        RECT 115.250 47.980 116.280 48.240 ;
        RECT 120.585 47.980 121.615 48.240 ;
        RECT 41.290 47.970 41.660 47.980 ;
        RECT 46.625 47.970 46.995 47.980 ;
        RECT 51.950 47.970 52.320 47.980 ;
        RECT 57.285 47.970 57.655 47.980 ;
        RECT 62.610 47.970 62.980 47.980 ;
        RECT 67.945 47.970 68.315 47.980 ;
        RECT 73.270 47.970 73.640 47.980 ;
        RECT 78.605 47.970 78.975 47.980 ;
        RECT 83.930 47.970 84.300 47.980 ;
        RECT 89.265 47.970 89.635 47.980 ;
        RECT 94.590 47.970 94.960 47.980 ;
        RECT 99.925 47.970 100.295 47.980 ;
        RECT 105.250 47.970 105.620 47.980 ;
        RECT 110.585 47.970 110.955 47.980 ;
        RECT 115.910 47.970 116.280 47.980 ;
        RECT 121.245 47.970 121.615 47.980 ;
        RECT 36.790 46.505 37.160 46.515 ;
        RECT 42.125 46.505 42.495 46.515 ;
        RECT 47.450 46.505 47.820 46.515 ;
        RECT 52.785 46.505 53.155 46.515 ;
        RECT 58.110 46.505 58.480 46.515 ;
        RECT 63.445 46.505 63.815 46.515 ;
        RECT 68.770 46.505 69.140 46.515 ;
        RECT 74.105 46.505 74.475 46.515 ;
        RECT 79.430 46.505 79.800 46.515 ;
        RECT 84.765 46.505 85.135 46.515 ;
        RECT 90.090 46.505 90.460 46.515 ;
        RECT 95.425 46.505 95.795 46.515 ;
        RECT 100.750 46.505 101.120 46.515 ;
        RECT 106.085 46.505 106.455 46.515 ;
        RECT 111.410 46.505 111.780 46.515 ;
        RECT 116.745 46.505 117.115 46.515 ;
        RECT 36.790 46.245 37.810 46.505 ;
        RECT 42.125 46.245 43.145 46.505 ;
        RECT 47.450 46.245 48.470 46.505 ;
        RECT 52.785 46.245 53.805 46.505 ;
        RECT 58.110 46.245 59.130 46.505 ;
        RECT 63.445 46.245 64.465 46.505 ;
        RECT 68.770 46.245 69.790 46.505 ;
        RECT 74.105 46.245 75.125 46.505 ;
        RECT 79.430 46.245 80.450 46.505 ;
        RECT 84.765 46.245 85.785 46.505 ;
        RECT 90.090 46.245 91.110 46.505 ;
        RECT 95.425 46.245 96.445 46.505 ;
        RECT 100.750 46.245 101.770 46.505 ;
        RECT 106.085 46.245 107.105 46.505 ;
        RECT 111.410 46.245 112.430 46.505 ;
        RECT 116.745 46.245 117.765 46.505 ;
        RECT 36.790 46.235 37.160 46.245 ;
        RECT 42.125 46.235 42.495 46.245 ;
        RECT 47.450 46.235 47.820 46.245 ;
        RECT 52.785 46.235 53.155 46.245 ;
        RECT 58.110 46.235 58.480 46.245 ;
        RECT 63.445 46.235 63.815 46.245 ;
        RECT 68.770 46.235 69.140 46.245 ;
        RECT 74.105 46.235 74.475 46.245 ;
        RECT 79.430 46.235 79.800 46.245 ;
        RECT 84.765 46.235 85.135 46.245 ;
        RECT 90.090 46.235 90.460 46.245 ;
        RECT 95.425 46.235 95.795 46.245 ;
        RECT 100.750 46.235 101.120 46.245 ;
        RECT 106.085 46.235 106.455 46.245 ;
        RECT 111.410 46.235 111.780 46.245 ;
        RECT 116.745 46.235 117.115 46.245 ;
        RECT 41.285 45.855 41.655 45.865 ;
        RECT 46.620 45.855 46.990 45.865 ;
        RECT 51.945 45.855 52.315 45.865 ;
        RECT 57.280 45.855 57.650 45.865 ;
        RECT 62.605 45.855 62.975 45.865 ;
        RECT 67.940 45.855 68.310 45.865 ;
        RECT 73.265 45.855 73.635 45.865 ;
        RECT 78.600 45.855 78.970 45.865 ;
        RECT 83.925 45.855 84.295 45.865 ;
        RECT 89.260 45.855 89.630 45.865 ;
        RECT 94.585 45.855 94.955 45.865 ;
        RECT 99.920 45.855 100.290 45.865 ;
        RECT 105.245 45.855 105.615 45.865 ;
        RECT 110.580 45.855 110.950 45.865 ;
        RECT 115.905 45.855 116.275 45.865 ;
        RECT 121.240 45.855 121.610 45.865 ;
        RECT 28.415 45.240 28.695 45.610 ;
        RECT 40.580 45.595 41.655 45.855 ;
        RECT 45.915 45.595 46.990 45.855 ;
        RECT 51.240 45.595 52.315 45.855 ;
        RECT 56.575 45.595 57.650 45.855 ;
        RECT 61.900 45.595 62.975 45.855 ;
        RECT 67.235 45.595 68.310 45.855 ;
        RECT 72.560 45.595 73.635 45.855 ;
        RECT 77.895 45.595 78.970 45.855 ;
        RECT 83.220 45.595 84.295 45.855 ;
        RECT 88.555 45.595 89.630 45.855 ;
        RECT 93.880 45.595 94.955 45.855 ;
        RECT 99.215 45.595 100.290 45.855 ;
        RECT 104.540 45.595 105.615 45.855 ;
        RECT 109.875 45.595 110.950 45.855 ;
        RECT 115.200 45.595 116.275 45.855 ;
        RECT 120.535 45.595 121.610 45.855 ;
        RECT 41.285 45.585 41.655 45.595 ;
        RECT 46.620 45.585 46.990 45.595 ;
        RECT 51.945 45.585 52.315 45.595 ;
        RECT 57.280 45.585 57.650 45.595 ;
        RECT 62.605 45.585 62.975 45.595 ;
        RECT 67.940 45.585 68.310 45.595 ;
        RECT 73.265 45.585 73.635 45.595 ;
        RECT 78.600 45.585 78.970 45.595 ;
        RECT 83.925 45.585 84.295 45.595 ;
        RECT 89.260 45.585 89.630 45.595 ;
        RECT 94.585 45.585 94.955 45.595 ;
        RECT 99.920 45.585 100.290 45.595 ;
        RECT 105.245 45.585 105.615 45.595 ;
        RECT 110.580 45.585 110.950 45.595 ;
        RECT 115.905 45.585 116.275 45.595 ;
        RECT 121.240 45.585 121.610 45.595 ;
        RECT 28.035 43.950 28.315 44.320 ;
        RECT 28.085 41.695 28.265 43.950 ;
        RECT 28.465 42.990 28.645 45.240 ;
        RECT 32.625 44.880 34.390 45.160 ;
        RECT 37.950 44.880 38.470 45.160 ;
        RECT 38.715 44.880 39.110 45.160 ;
        RECT 39.330 44.880 39.730 45.160 ;
        RECT 43.285 44.880 43.805 45.160 ;
        RECT 44.050 44.880 44.445 45.160 ;
        RECT 44.665 44.880 45.065 45.160 ;
        RECT 48.610 44.880 49.130 45.160 ;
        RECT 49.375 44.880 49.770 45.160 ;
        RECT 49.990 44.880 50.390 45.160 ;
        RECT 53.945 44.880 54.465 45.160 ;
        RECT 54.710 44.880 55.105 45.160 ;
        RECT 55.325 44.880 55.725 45.160 ;
        RECT 59.270 44.880 59.790 45.160 ;
        RECT 60.035 44.880 60.430 45.160 ;
        RECT 60.650 44.880 61.050 45.160 ;
        RECT 64.605 44.880 65.125 45.160 ;
        RECT 65.370 44.880 65.765 45.160 ;
        RECT 65.985 44.880 66.385 45.160 ;
        RECT 69.930 44.880 70.450 45.160 ;
        RECT 70.695 44.880 71.090 45.160 ;
        RECT 71.310 44.880 71.710 45.160 ;
        RECT 75.265 44.880 75.785 45.160 ;
        RECT 76.030 44.880 76.425 45.160 ;
        RECT 76.645 44.880 77.045 45.160 ;
        RECT 80.590 44.880 81.110 45.160 ;
        RECT 81.355 44.880 81.750 45.160 ;
        RECT 81.970 44.880 82.370 45.160 ;
        RECT 85.925 44.880 86.445 45.160 ;
        RECT 86.690 44.880 87.085 45.160 ;
        RECT 87.305 44.880 87.705 45.160 ;
        RECT 91.250 44.880 91.770 45.160 ;
        RECT 92.015 44.880 92.410 45.160 ;
        RECT 92.630 44.880 93.030 45.160 ;
        RECT 96.585 44.880 97.105 45.160 ;
        RECT 97.350 44.880 97.745 45.160 ;
        RECT 97.965 44.880 98.365 45.160 ;
        RECT 101.910 44.880 102.430 45.160 ;
        RECT 102.675 44.880 103.070 45.160 ;
        RECT 103.290 44.880 103.690 45.160 ;
        RECT 107.245 44.880 107.765 45.160 ;
        RECT 108.010 44.880 108.405 45.160 ;
        RECT 108.625 44.880 109.025 45.160 ;
        RECT 112.570 44.880 113.090 45.160 ;
        RECT 113.335 44.880 113.730 45.160 ;
        RECT 113.950 44.880 114.350 45.160 ;
        RECT 117.905 44.880 118.425 45.160 ;
        RECT 118.670 44.880 119.065 45.160 ;
        RECT 119.285 44.880 119.685 45.160 ;
        RECT 123.230 44.880 124.995 45.160 ;
        RECT 36.785 44.660 37.155 44.670 ;
        RECT 42.120 44.660 42.490 44.670 ;
        RECT 47.445 44.660 47.815 44.670 ;
        RECT 52.780 44.660 53.150 44.670 ;
        RECT 58.105 44.660 58.475 44.670 ;
        RECT 63.440 44.660 63.810 44.670 ;
        RECT 68.765 44.660 69.135 44.670 ;
        RECT 74.100 44.660 74.470 44.670 ;
        RECT 79.425 44.660 79.795 44.670 ;
        RECT 84.760 44.660 85.130 44.670 ;
        RECT 90.085 44.660 90.455 44.670 ;
        RECT 95.420 44.660 95.790 44.670 ;
        RECT 100.745 44.660 101.115 44.670 ;
        RECT 106.080 44.660 106.450 44.670 ;
        RECT 111.405 44.660 111.775 44.670 ;
        RECT 116.740 44.660 117.110 44.670 ;
        RECT 36.785 44.400 37.810 44.660 ;
        RECT 41.285 44.570 41.655 44.580 ;
        RECT 36.785 44.390 37.155 44.400 ;
        RECT 40.630 44.310 41.655 44.570 ;
        RECT 42.120 44.400 43.145 44.660 ;
        RECT 46.620 44.570 46.990 44.580 ;
        RECT 42.120 44.390 42.490 44.400 ;
        RECT 45.965 44.310 46.990 44.570 ;
        RECT 47.445 44.400 48.470 44.660 ;
        RECT 51.945 44.570 52.315 44.580 ;
        RECT 47.445 44.390 47.815 44.400 ;
        RECT 51.290 44.310 52.315 44.570 ;
        RECT 52.780 44.400 53.805 44.660 ;
        RECT 57.280 44.570 57.650 44.580 ;
        RECT 52.780 44.390 53.150 44.400 ;
        RECT 56.625 44.310 57.650 44.570 ;
        RECT 58.105 44.400 59.130 44.660 ;
        RECT 62.605 44.570 62.975 44.580 ;
        RECT 58.105 44.390 58.475 44.400 ;
        RECT 61.950 44.310 62.975 44.570 ;
        RECT 63.440 44.400 64.465 44.660 ;
        RECT 67.940 44.570 68.310 44.580 ;
        RECT 63.440 44.390 63.810 44.400 ;
        RECT 67.285 44.310 68.310 44.570 ;
        RECT 68.765 44.400 69.790 44.660 ;
        RECT 73.265 44.570 73.635 44.580 ;
        RECT 68.765 44.390 69.135 44.400 ;
        RECT 72.610 44.310 73.635 44.570 ;
        RECT 74.100 44.400 75.125 44.660 ;
        RECT 78.600 44.570 78.970 44.580 ;
        RECT 74.100 44.390 74.470 44.400 ;
        RECT 77.945 44.310 78.970 44.570 ;
        RECT 79.425 44.400 80.450 44.660 ;
        RECT 83.925 44.570 84.295 44.580 ;
        RECT 79.425 44.390 79.795 44.400 ;
        RECT 83.270 44.310 84.295 44.570 ;
        RECT 84.760 44.400 85.785 44.660 ;
        RECT 89.260 44.570 89.630 44.580 ;
        RECT 84.760 44.390 85.130 44.400 ;
        RECT 88.605 44.310 89.630 44.570 ;
        RECT 90.085 44.400 91.110 44.660 ;
        RECT 94.585 44.570 94.955 44.580 ;
        RECT 90.085 44.390 90.455 44.400 ;
        RECT 93.930 44.310 94.955 44.570 ;
        RECT 95.420 44.400 96.445 44.660 ;
        RECT 99.920 44.570 100.290 44.580 ;
        RECT 95.420 44.390 95.790 44.400 ;
        RECT 99.265 44.310 100.290 44.570 ;
        RECT 100.745 44.400 101.770 44.660 ;
        RECT 105.245 44.570 105.615 44.580 ;
        RECT 100.745 44.390 101.115 44.400 ;
        RECT 104.590 44.310 105.615 44.570 ;
        RECT 106.080 44.400 107.105 44.660 ;
        RECT 110.580 44.570 110.950 44.580 ;
        RECT 106.080 44.390 106.450 44.400 ;
        RECT 109.925 44.310 110.950 44.570 ;
        RECT 111.405 44.400 112.430 44.660 ;
        RECT 115.905 44.570 116.275 44.580 ;
        RECT 111.405 44.390 111.775 44.400 ;
        RECT 115.250 44.310 116.275 44.570 ;
        RECT 116.740 44.400 117.765 44.660 ;
        RECT 121.240 44.570 121.610 44.580 ;
        RECT 116.740 44.390 117.110 44.400 ;
        RECT 120.585 44.310 121.610 44.570 ;
        RECT 41.285 44.300 41.655 44.310 ;
        RECT 46.620 44.300 46.990 44.310 ;
        RECT 51.945 44.300 52.315 44.310 ;
        RECT 57.280 44.300 57.650 44.310 ;
        RECT 62.605 44.300 62.975 44.310 ;
        RECT 67.940 44.300 68.310 44.310 ;
        RECT 73.265 44.300 73.635 44.310 ;
        RECT 78.600 44.300 78.970 44.310 ;
        RECT 83.925 44.300 84.295 44.310 ;
        RECT 89.260 44.300 89.630 44.310 ;
        RECT 94.585 44.300 94.955 44.310 ;
        RECT 99.920 44.300 100.290 44.310 ;
        RECT 105.245 44.300 105.615 44.310 ;
        RECT 110.580 44.300 110.950 44.310 ;
        RECT 115.905 44.300 116.275 44.310 ;
        RECT 121.240 44.300 121.610 44.310 ;
        RECT 28.410 42.620 28.690 42.990 ;
        RECT 36.785 42.635 37.155 42.645 ;
        RECT 42.120 42.635 42.490 42.645 ;
        RECT 47.445 42.635 47.815 42.645 ;
        RECT 52.780 42.635 53.150 42.645 ;
        RECT 58.105 42.635 58.475 42.645 ;
        RECT 63.440 42.635 63.810 42.645 ;
        RECT 68.765 42.635 69.135 42.645 ;
        RECT 74.100 42.635 74.470 42.645 ;
        RECT 79.425 42.635 79.795 42.645 ;
        RECT 84.760 42.635 85.130 42.645 ;
        RECT 90.085 42.635 90.455 42.645 ;
        RECT 95.420 42.635 95.790 42.645 ;
        RECT 100.745 42.635 101.115 42.645 ;
        RECT 106.080 42.635 106.450 42.645 ;
        RECT 111.405 42.635 111.775 42.645 ;
        RECT 116.740 42.635 117.110 42.645 ;
        RECT 28.035 41.325 28.315 41.695 ;
        RECT 28.085 38.075 28.265 41.325 ;
        RECT 28.035 37.705 28.315 38.075 ;
        RECT 28.085 35.455 28.265 37.705 ;
        RECT 28.465 36.785 28.645 42.620 ;
        RECT 36.785 42.375 37.810 42.635 ;
        RECT 41.285 42.540 41.655 42.550 ;
        RECT 36.785 42.365 37.155 42.375 ;
        RECT 40.630 42.280 41.655 42.540 ;
        RECT 42.120 42.375 43.145 42.635 ;
        RECT 46.620 42.540 46.990 42.550 ;
        RECT 42.120 42.365 42.490 42.375 ;
        RECT 45.965 42.280 46.990 42.540 ;
        RECT 47.445 42.375 48.470 42.635 ;
        RECT 51.945 42.540 52.315 42.550 ;
        RECT 47.445 42.365 47.815 42.375 ;
        RECT 51.290 42.280 52.315 42.540 ;
        RECT 52.780 42.375 53.805 42.635 ;
        RECT 57.280 42.540 57.650 42.550 ;
        RECT 52.780 42.365 53.150 42.375 ;
        RECT 56.625 42.280 57.650 42.540 ;
        RECT 58.105 42.375 59.130 42.635 ;
        RECT 62.605 42.540 62.975 42.550 ;
        RECT 58.105 42.365 58.475 42.375 ;
        RECT 61.950 42.280 62.975 42.540 ;
        RECT 63.440 42.375 64.465 42.635 ;
        RECT 67.940 42.540 68.310 42.550 ;
        RECT 63.440 42.365 63.810 42.375 ;
        RECT 67.285 42.280 68.310 42.540 ;
        RECT 68.765 42.375 69.790 42.635 ;
        RECT 73.265 42.540 73.635 42.550 ;
        RECT 68.765 42.365 69.135 42.375 ;
        RECT 72.610 42.280 73.635 42.540 ;
        RECT 74.100 42.375 75.125 42.635 ;
        RECT 78.600 42.540 78.970 42.550 ;
        RECT 74.100 42.365 74.470 42.375 ;
        RECT 77.945 42.280 78.970 42.540 ;
        RECT 79.425 42.375 80.450 42.635 ;
        RECT 83.925 42.540 84.295 42.550 ;
        RECT 79.425 42.365 79.795 42.375 ;
        RECT 83.270 42.280 84.295 42.540 ;
        RECT 84.760 42.375 85.785 42.635 ;
        RECT 89.260 42.540 89.630 42.550 ;
        RECT 84.760 42.365 85.130 42.375 ;
        RECT 88.605 42.280 89.630 42.540 ;
        RECT 90.085 42.375 91.110 42.635 ;
        RECT 94.585 42.540 94.955 42.550 ;
        RECT 90.085 42.365 90.455 42.375 ;
        RECT 93.930 42.280 94.955 42.540 ;
        RECT 95.420 42.375 96.445 42.635 ;
        RECT 99.920 42.540 100.290 42.550 ;
        RECT 95.420 42.365 95.790 42.375 ;
        RECT 99.265 42.280 100.290 42.540 ;
        RECT 100.745 42.375 101.770 42.635 ;
        RECT 105.245 42.540 105.615 42.550 ;
        RECT 100.745 42.365 101.115 42.375 ;
        RECT 104.590 42.280 105.615 42.540 ;
        RECT 106.080 42.375 107.105 42.635 ;
        RECT 110.580 42.540 110.950 42.550 ;
        RECT 106.080 42.365 106.450 42.375 ;
        RECT 109.925 42.280 110.950 42.540 ;
        RECT 111.405 42.375 112.430 42.635 ;
        RECT 115.905 42.540 116.275 42.550 ;
        RECT 111.405 42.365 111.775 42.375 ;
        RECT 115.250 42.280 116.275 42.540 ;
        RECT 116.740 42.375 117.765 42.635 ;
        RECT 121.240 42.540 121.610 42.550 ;
        RECT 116.740 42.365 117.110 42.375 ;
        RECT 120.585 42.280 121.610 42.540 ;
        RECT 41.285 42.270 41.655 42.280 ;
        RECT 46.620 42.270 46.990 42.280 ;
        RECT 51.945 42.270 52.315 42.280 ;
        RECT 57.280 42.270 57.650 42.280 ;
        RECT 62.605 42.270 62.975 42.280 ;
        RECT 67.940 42.270 68.310 42.280 ;
        RECT 73.265 42.270 73.635 42.280 ;
        RECT 78.600 42.270 78.970 42.280 ;
        RECT 83.925 42.270 84.295 42.280 ;
        RECT 89.260 42.270 89.630 42.280 ;
        RECT 94.585 42.270 94.955 42.280 ;
        RECT 99.920 42.270 100.290 42.280 ;
        RECT 105.245 42.270 105.615 42.280 ;
        RECT 110.580 42.270 110.950 42.280 ;
        RECT 115.905 42.270 116.275 42.280 ;
        RECT 121.240 42.270 121.610 42.280 ;
        RECT 34.005 41.985 34.400 41.990 ;
        RECT 33.390 41.705 35.160 41.985 ;
        RECT 38.715 41.705 39.110 41.985 ;
        RECT 39.330 41.710 39.755 41.990 ;
        RECT 40.120 41.705 41.015 41.985 ;
        RECT 44.050 41.705 44.445 41.985 ;
        RECT 44.665 41.710 45.090 41.990 ;
        RECT 45.455 41.705 46.350 41.985 ;
        RECT 49.375 41.705 49.770 41.985 ;
        RECT 49.990 41.710 50.415 41.990 ;
        RECT 50.780 41.705 51.675 41.985 ;
        RECT 54.710 41.705 55.105 41.985 ;
        RECT 55.325 41.710 55.750 41.990 ;
        RECT 56.115 41.705 57.010 41.985 ;
        RECT 60.035 41.705 60.430 41.985 ;
        RECT 60.650 41.710 61.075 41.990 ;
        RECT 61.440 41.705 62.335 41.985 ;
        RECT 65.370 41.705 65.765 41.985 ;
        RECT 65.985 41.710 66.410 41.990 ;
        RECT 66.775 41.705 67.670 41.985 ;
        RECT 70.695 41.705 71.090 41.985 ;
        RECT 71.310 41.710 71.735 41.990 ;
        RECT 72.100 41.705 72.995 41.985 ;
        RECT 76.030 41.705 76.425 41.985 ;
        RECT 76.645 41.710 77.070 41.990 ;
        RECT 77.435 41.705 78.330 41.985 ;
        RECT 81.355 41.705 81.750 41.985 ;
        RECT 81.970 41.710 82.395 41.990 ;
        RECT 82.760 41.705 83.655 41.985 ;
        RECT 86.690 41.705 87.085 41.985 ;
        RECT 87.305 41.710 87.730 41.990 ;
        RECT 88.095 41.705 88.990 41.985 ;
        RECT 92.015 41.705 92.410 41.985 ;
        RECT 92.630 41.710 93.055 41.990 ;
        RECT 93.420 41.705 94.315 41.985 ;
        RECT 97.350 41.705 97.745 41.985 ;
        RECT 97.965 41.710 98.390 41.990 ;
        RECT 98.755 41.705 99.650 41.985 ;
        RECT 102.675 41.705 103.070 41.985 ;
        RECT 103.290 41.710 103.715 41.990 ;
        RECT 104.080 41.705 104.975 41.985 ;
        RECT 108.010 41.705 108.405 41.985 ;
        RECT 108.625 41.710 109.050 41.990 ;
        RECT 109.415 41.705 110.310 41.985 ;
        RECT 113.335 41.705 113.730 41.985 ;
        RECT 113.950 41.710 114.375 41.990 ;
        RECT 114.740 41.705 115.635 41.985 ;
        RECT 118.670 41.705 119.065 41.985 ;
        RECT 119.285 41.710 119.710 41.990 ;
        RECT 124.610 41.985 125.005 41.990 ;
        RECT 120.075 41.705 120.970 41.985 ;
        RECT 123.995 41.705 125.765 41.985 ;
        RECT 36.785 41.335 37.155 41.345 ;
        RECT 42.120 41.335 42.490 41.345 ;
        RECT 47.445 41.335 47.815 41.345 ;
        RECT 52.780 41.335 53.150 41.345 ;
        RECT 58.105 41.335 58.475 41.345 ;
        RECT 63.440 41.335 63.810 41.345 ;
        RECT 68.765 41.335 69.135 41.345 ;
        RECT 74.100 41.335 74.470 41.345 ;
        RECT 79.425 41.335 79.795 41.345 ;
        RECT 84.760 41.335 85.130 41.345 ;
        RECT 90.085 41.335 90.455 41.345 ;
        RECT 95.420 41.335 95.790 41.345 ;
        RECT 100.745 41.335 101.115 41.345 ;
        RECT 106.080 41.335 106.450 41.345 ;
        RECT 111.405 41.335 111.775 41.345 ;
        RECT 116.740 41.335 117.110 41.345 ;
        RECT 36.785 41.075 37.860 41.335 ;
        RECT 42.120 41.075 43.195 41.335 ;
        RECT 47.445 41.075 48.520 41.335 ;
        RECT 52.780 41.075 53.855 41.335 ;
        RECT 58.105 41.075 59.180 41.335 ;
        RECT 63.440 41.075 64.515 41.335 ;
        RECT 68.765 41.075 69.840 41.335 ;
        RECT 74.100 41.075 75.175 41.335 ;
        RECT 79.425 41.075 80.500 41.335 ;
        RECT 84.760 41.075 85.835 41.335 ;
        RECT 90.085 41.075 91.160 41.335 ;
        RECT 95.420 41.075 96.495 41.335 ;
        RECT 100.745 41.075 101.820 41.335 ;
        RECT 106.080 41.075 107.155 41.335 ;
        RECT 111.405 41.075 112.480 41.335 ;
        RECT 116.740 41.075 117.815 41.335 ;
        RECT 36.785 41.065 37.155 41.075 ;
        RECT 42.120 41.065 42.490 41.075 ;
        RECT 47.445 41.065 47.815 41.075 ;
        RECT 52.780 41.065 53.150 41.075 ;
        RECT 58.105 41.065 58.475 41.075 ;
        RECT 63.440 41.065 63.810 41.075 ;
        RECT 68.765 41.065 69.135 41.075 ;
        RECT 74.100 41.065 74.470 41.075 ;
        RECT 79.425 41.065 79.795 41.075 ;
        RECT 84.760 41.065 85.130 41.075 ;
        RECT 90.085 41.065 90.455 41.075 ;
        RECT 95.420 41.065 95.790 41.075 ;
        RECT 100.745 41.065 101.115 41.075 ;
        RECT 106.080 41.065 106.450 41.075 ;
        RECT 111.405 41.065 111.775 41.075 ;
        RECT 116.740 41.065 117.110 41.075 ;
        RECT 41.290 40.705 41.660 40.715 ;
        RECT 46.625 40.705 46.995 40.715 ;
        RECT 51.950 40.705 52.320 40.715 ;
        RECT 57.285 40.705 57.655 40.715 ;
        RECT 62.610 40.705 62.980 40.715 ;
        RECT 67.945 40.705 68.315 40.715 ;
        RECT 73.270 40.705 73.640 40.715 ;
        RECT 78.605 40.705 78.975 40.715 ;
        RECT 83.930 40.705 84.300 40.715 ;
        RECT 89.265 40.705 89.635 40.715 ;
        RECT 94.590 40.705 94.960 40.715 ;
        RECT 99.925 40.705 100.295 40.715 ;
        RECT 105.250 40.705 105.620 40.715 ;
        RECT 110.585 40.705 110.955 40.715 ;
        RECT 115.910 40.705 116.280 40.715 ;
        RECT 121.245 40.705 121.615 40.715 ;
        RECT 40.630 40.445 41.660 40.705 ;
        RECT 45.965 40.445 46.995 40.705 ;
        RECT 51.290 40.445 52.320 40.705 ;
        RECT 56.625 40.445 57.655 40.705 ;
        RECT 61.950 40.445 62.980 40.705 ;
        RECT 67.285 40.445 68.315 40.705 ;
        RECT 72.610 40.445 73.640 40.705 ;
        RECT 77.945 40.445 78.975 40.705 ;
        RECT 83.270 40.445 84.300 40.705 ;
        RECT 88.605 40.445 89.635 40.705 ;
        RECT 93.930 40.445 94.960 40.705 ;
        RECT 99.265 40.445 100.295 40.705 ;
        RECT 104.590 40.445 105.620 40.705 ;
        RECT 109.925 40.445 110.955 40.705 ;
        RECT 115.250 40.445 116.280 40.705 ;
        RECT 120.585 40.445 121.615 40.705 ;
        RECT 41.290 40.435 41.660 40.445 ;
        RECT 46.625 40.435 46.995 40.445 ;
        RECT 51.950 40.435 52.320 40.445 ;
        RECT 57.285 40.435 57.655 40.445 ;
        RECT 62.610 40.435 62.980 40.445 ;
        RECT 67.945 40.435 68.315 40.445 ;
        RECT 73.270 40.435 73.640 40.445 ;
        RECT 78.605 40.435 78.975 40.445 ;
        RECT 83.930 40.435 84.300 40.445 ;
        RECT 89.265 40.435 89.635 40.445 ;
        RECT 94.590 40.435 94.960 40.445 ;
        RECT 99.925 40.435 100.295 40.445 ;
        RECT 105.250 40.435 105.620 40.445 ;
        RECT 110.585 40.435 110.955 40.445 ;
        RECT 115.910 40.435 116.280 40.445 ;
        RECT 121.245 40.435 121.615 40.445 ;
        RECT 36.790 38.970 37.160 38.980 ;
        RECT 42.125 38.970 42.495 38.980 ;
        RECT 47.450 38.970 47.820 38.980 ;
        RECT 52.785 38.970 53.155 38.980 ;
        RECT 58.110 38.970 58.480 38.980 ;
        RECT 63.445 38.970 63.815 38.980 ;
        RECT 68.770 38.970 69.140 38.980 ;
        RECT 74.105 38.970 74.475 38.980 ;
        RECT 79.430 38.970 79.800 38.980 ;
        RECT 84.765 38.970 85.135 38.980 ;
        RECT 90.090 38.970 90.460 38.980 ;
        RECT 95.425 38.970 95.795 38.980 ;
        RECT 100.750 38.970 101.120 38.980 ;
        RECT 106.085 38.970 106.455 38.980 ;
        RECT 111.410 38.970 111.780 38.980 ;
        RECT 116.745 38.970 117.115 38.980 ;
        RECT 36.790 38.710 37.810 38.970 ;
        RECT 42.125 38.710 43.145 38.970 ;
        RECT 47.450 38.710 48.470 38.970 ;
        RECT 52.785 38.710 53.805 38.970 ;
        RECT 58.110 38.710 59.130 38.970 ;
        RECT 63.445 38.710 64.465 38.970 ;
        RECT 68.770 38.710 69.790 38.970 ;
        RECT 74.105 38.710 75.125 38.970 ;
        RECT 79.430 38.710 80.450 38.970 ;
        RECT 84.765 38.710 85.785 38.970 ;
        RECT 90.090 38.710 91.110 38.970 ;
        RECT 95.425 38.710 96.445 38.970 ;
        RECT 100.750 38.710 101.770 38.970 ;
        RECT 106.085 38.710 107.105 38.970 ;
        RECT 111.410 38.710 112.430 38.970 ;
        RECT 116.745 38.710 117.765 38.970 ;
        RECT 36.790 38.700 37.160 38.710 ;
        RECT 42.125 38.700 42.495 38.710 ;
        RECT 47.450 38.700 47.820 38.710 ;
        RECT 52.785 38.700 53.155 38.710 ;
        RECT 58.110 38.700 58.480 38.710 ;
        RECT 63.445 38.700 63.815 38.710 ;
        RECT 68.770 38.700 69.140 38.710 ;
        RECT 74.105 38.700 74.475 38.710 ;
        RECT 79.430 38.700 79.800 38.710 ;
        RECT 84.765 38.700 85.135 38.710 ;
        RECT 90.090 38.700 90.460 38.710 ;
        RECT 95.425 38.700 95.795 38.710 ;
        RECT 100.750 38.700 101.120 38.710 ;
        RECT 106.085 38.700 106.455 38.710 ;
        RECT 111.410 38.700 111.780 38.710 ;
        RECT 116.745 38.700 117.115 38.710 ;
        RECT 41.285 38.320 41.655 38.330 ;
        RECT 46.620 38.320 46.990 38.330 ;
        RECT 51.945 38.320 52.315 38.330 ;
        RECT 57.280 38.320 57.650 38.330 ;
        RECT 62.605 38.320 62.975 38.330 ;
        RECT 67.940 38.320 68.310 38.330 ;
        RECT 73.265 38.320 73.635 38.330 ;
        RECT 78.600 38.320 78.970 38.330 ;
        RECT 83.925 38.320 84.295 38.330 ;
        RECT 89.260 38.320 89.630 38.330 ;
        RECT 94.585 38.320 94.955 38.330 ;
        RECT 99.920 38.320 100.290 38.330 ;
        RECT 105.245 38.320 105.615 38.330 ;
        RECT 110.580 38.320 110.950 38.330 ;
        RECT 115.905 38.320 116.275 38.330 ;
        RECT 121.240 38.320 121.610 38.330 ;
        RECT 40.580 38.060 41.655 38.320 ;
        RECT 45.915 38.060 46.990 38.320 ;
        RECT 51.240 38.060 52.315 38.320 ;
        RECT 56.575 38.060 57.650 38.320 ;
        RECT 61.900 38.060 62.975 38.320 ;
        RECT 67.235 38.060 68.310 38.320 ;
        RECT 72.560 38.060 73.635 38.320 ;
        RECT 77.895 38.060 78.970 38.320 ;
        RECT 83.220 38.060 84.295 38.320 ;
        RECT 88.555 38.060 89.630 38.320 ;
        RECT 93.880 38.060 94.955 38.320 ;
        RECT 99.215 38.060 100.290 38.320 ;
        RECT 104.540 38.060 105.615 38.320 ;
        RECT 109.875 38.060 110.950 38.320 ;
        RECT 115.200 38.060 116.275 38.320 ;
        RECT 120.535 38.060 121.610 38.320 ;
        RECT 41.285 38.050 41.655 38.060 ;
        RECT 46.620 38.050 46.990 38.060 ;
        RECT 51.945 38.050 52.315 38.060 ;
        RECT 57.280 38.050 57.650 38.060 ;
        RECT 62.605 38.050 62.975 38.060 ;
        RECT 67.940 38.050 68.310 38.060 ;
        RECT 73.265 38.050 73.635 38.060 ;
        RECT 78.600 38.050 78.970 38.060 ;
        RECT 83.925 38.050 84.295 38.060 ;
        RECT 89.260 38.050 89.630 38.060 ;
        RECT 94.585 38.050 94.955 38.060 ;
        RECT 99.920 38.050 100.290 38.060 ;
        RECT 105.245 38.050 105.615 38.060 ;
        RECT 110.580 38.050 110.950 38.060 ;
        RECT 115.905 38.050 116.275 38.060 ;
        RECT 121.240 38.050 121.610 38.060 ;
        RECT 32.625 37.345 34.390 37.625 ;
        RECT 37.430 37.345 38.320 37.625 ;
        RECT 38.715 37.345 39.110 37.625 ;
        RECT 39.330 37.345 39.715 37.625 ;
        RECT 42.765 37.345 43.655 37.625 ;
        RECT 44.050 37.345 44.445 37.625 ;
        RECT 44.665 37.345 45.050 37.625 ;
        RECT 48.090 37.345 48.980 37.625 ;
        RECT 49.375 37.345 49.770 37.625 ;
        RECT 49.990 37.345 50.375 37.625 ;
        RECT 53.425 37.345 54.315 37.625 ;
        RECT 54.710 37.345 55.105 37.625 ;
        RECT 55.325 37.345 55.710 37.625 ;
        RECT 58.750 37.345 59.640 37.625 ;
        RECT 60.035 37.345 60.430 37.625 ;
        RECT 60.650 37.345 61.035 37.625 ;
        RECT 64.085 37.345 64.975 37.625 ;
        RECT 65.370 37.345 65.765 37.625 ;
        RECT 65.985 37.345 66.370 37.625 ;
        RECT 69.410 37.345 70.300 37.625 ;
        RECT 70.695 37.345 71.090 37.625 ;
        RECT 71.310 37.345 71.695 37.625 ;
        RECT 74.745 37.345 75.635 37.625 ;
        RECT 76.030 37.345 76.425 37.625 ;
        RECT 76.645 37.345 77.030 37.625 ;
        RECT 80.070 37.345 80.960 37.625 ;
        RECT 81.355 37.345 81.750 37.625 ;
        RECT 81.970 37.345 82.355 37.625 ;
        RECT 85.405 37.345 86.295 37.625 ;
        RECT 86.690 37.345 87.085 37.625 ;
        RECT 87.305 37.345 87.690 37.625 ;
        RECT 90.730 37.345 91.620 37.625 ;
        RECT 92.015 37.345 92.410 37.625 ;
        RECT 92.630 37.345 93.015 37.625 ;
        RECT 96.065 37.345 96.955 37.625 ;
        RECT 97.350 37.345 97.745 37.625 ;
        RECT 97.965 37.345 98.350 37.625 ;
        RECT 101.390 37.345 102.280 37.625 ;
        RECT 102.675 37.345 103.070 37.625 ;
        RECT 103.290 37.345 103.675 37.625 ;
        RECT 106.725 37.345 107.615 37.625 ;
        RECT 108.010 37.345 108.405 37.625 ;
        RECT 108.625 37.345 109.010 37.625 ;
        RECT 112.050 37.345 112.940 37.625 ;
        RECT 113.335 37.345 113.730 37.625 ;
        RECT 113.950 37.345 114.335 37.625 ;
        RECT 117.385 37.345 118.275 37.625 ;
        RECT 118.670 37.345 119.065 37.625 ;
        RECT 119.285 37.345 119.670 37.625 ;
        RECT 123.230 37.345 124.995 37.625 ;
        RECT 36.785 37.125 37.155 37.135 ;
        RECT 36.785 36.865 37.810 37.125 ;
        RECT 39.375 37.120 39.655 37.345 ;
        RECT 36.785 36.855 37.155 36.865 ;
        RECT 38.105 36.840 39.655 37.120 ;
        RECT 42.120 37.125 42.490 37.135 ;
        RECT 41.285 37.035 41.655 37.045 ;
        RECT 28.415 36.415 28.695 36.785 ;
        RECT 40.630 36.775 41.655 37.035 ;
        RECT 42.120 36.865 43.145 37.125 ;
        RECT 44.710 37.120 44.990 37.345 ;
        RECT 42.120 36.855 42.490 36.865 ;
        RECT 43.440 36.840 44.990 37.120 ;
        RECT 47.445 37.125 47.815 37.135 ;
        RECT 46.620 37.035 46.990 37.045 ;
        RECT 45.965 36.775 46.990 37.035 ;
        RECT 47.445 36.865 48.470 37.125 ;
        RECT 50.035 37.120 50.315 37.345 ;
        RECT 47.445 36.855 47.815 36.865 ;
        RECT 48.765 36.840 50.315 37.120 ;
        RECT 52.780 37.125 53.150 37.135 ;
        RECT 51.945 37.035 52.315 37.045 ;
        RECT 51.290 36.775 52.315 37.035 ;
        RECT 52.780 36.865 53.805 37.125 ;
        RECT 55.370 37.120 55.650 37.345 ;
        RECT 52.780 36.855 53.150 36.865 ;
        RECT 54.100 36.840 55.650 37.120 ;
        RECT 58.105 37.125 58.475 37.135 ;
        RECT 57.280 37.035 57.650 37.045 ;
        RECT 56.625 36.775 57.650 37.035 ;
        RECT 58.105 36.865 59.130 37.125 ;
        RECT 60.695 37.120 60.975 37.345 ;
        RECT 58.105 36.855 58.475 36.865 ;
        RECT 59.425 36.840 60.975 37.120 ;
        RECT 63.440 37.125 63.810 37.135 ;
        RECT 62.605 37.035 62.975 37.045 ;
        RECT 61.950 36.775 62.975 37.035 ;
        RECT 63.440 36.865 64.465 37.125 ;
        RECT 66.030 37.120 66.310 37.345 ;
        RECT 63.440 36.855 63.810 36.865 ;
        RECT 64.760 36.840 66.310 37.120 ;
        RECT 68.765 37.125 69.135 37.135 ;
        RECT 67.940 37.035 68.310 37.045 ;
        RECT 67.285 36.775 68.310 37.035 ;
        RECT 68.765 36.865 69.790 37.125 ;
        RECT 71.355 37.120 71.635 37.345 ;
        RECT 68.765 36.855 69.135 36.865 ;
        RECT 70.085 36.840 71.635 37.120 ;
        RECT 74.100 37.125 74.470 37.135 ;
        RECT 73.265 37.035 73.635 37.045 ;
        RECT 72.610 36.775 73.635 37.035 ;
        RECT 74.100 36.865 75.125 37.125 ;
        RECT 76.690 37.120 76.970 37.345 ;
        RECT 74.100 36.855 74.470 36.865 ;
        RECT 75.420 36.840 76.970 37.120 ;
        RECT 79.425 37.125 79.795 37.135 ;
        RECT 78.600 37.035 78.970 37.045 ;
        RECT 77.945 36.775 78.970 37.035 ;
        RECT 79.425 36.865 80.450 37.125 ;
        RECT 82.015 37.120 82.295 37.345 ;
        RECT 79.425 36.855 79.795 36.865 ;
        RECT 80.745 36.840 82.295 37.120 ;
        RECT 84.760 37.125 85.130 37.135 ;
        RECT 83.925 37.035 84.295 37.045 ;
        RECT 83.270 36.775 84.295 37.035 ;
        RECT 84.760 36.865 85.785 37.125 ;
        RECT 87.350 37.120 87.630 37.345 ;
        RECT 84.760 36.855 85.130 36.865 ;
        RECT 86.080 36.840 87.630 37.120 ;
        RECT 90.085 37.125 90.455 37.135 ;
        RECT 89.260 37.035 89.630 37.045 ;
        RECT 88.605 36.775 89.630 37.035 ;
        RECT 90.085 36.865 91.110 37.125 ;
        RECT 92.675 37.120 92.955 37.345 ;
        RECT 90.085 36.855 90.455 36.865 ;
        RECT 91.405 36.840 92.955 37.120 ;
        RECT 95.420 37.125 95.790 37.135 ;
        RECT 94.585 37.035 94.955 37.045 ;
        RECT 93.930 36.775 94.955 37.035 ;
        RECT 95.420 36.865 96.445 37.125 ;
        RECT 98.010 37.120 98.290 37.345 ;
        RECT 95.420 36.855 95.790 36.865 ;
        RECT 96.740 36.840 98.290 37.120 ;
        RECT 100.745 37.125 101.115 37.135 ;
        RECT 99.920 37.035 100.290 37.045 ;
        RECT 99.265 36.775 100.290 37.035 ;
        RECT 100.745 36.865 101.770 37.125 ;
        RECT 103.335 37.120 103.615 37.345 ;
        RECT 100.745 36.855 101.115 36.865 ;
        RECT 102.065 36.840 103.615 37.120 ;
        RECT 106.080 37.125 106.450 37.135 ;
        RECT 105.245 37.035 105.615 37.045 ;
        RECT 104.590 36.775 105.615 37.035 ;
        RECT 106.080 36.865 107.105 37.125 ;
        RECT 108.670 37.120 108.950 37.345 ;
        RECT 106.080 36.855 106.450 36.865 ;
        RECT 107.400 36.840 108.950 37.120 ;
        RECT 111.405 37.125 111.775 37.135 ;
        RECT 110.580 37.035 110.950 37.045 ;
        RECT 109.925 36.775 110.950 37.035 ;
        RECT 111.405 36.865 112.430 37.125 ;
        RECT 113.995 37.120 114.275 37.345 ;
        RECT 111.405 36.855 111.775 36.865 ;
        RECT 112.725 36.840 114.275 37.120 ;
        RECT 116.740 37.125 117.110 37.135 ;
        RECT 115.905 37.035 116.275 37.045 ;
        RECT 115.250 36.775 116.275 37.035 ;
        RECT 116.740 36.865 117.765 37.125 ;
        RECT 119.330 37.120 119.610 37.345 ;
        RECT 116.740 36.855 117.110 36.865 ;
        RECT 118.060 36.840 119.610 37.120 ;
        RECT 121.240 37.035 121.610 37.045 ;
        RECT 120.585 36.775 121.610 37.035 ;
        RECT 41.285 36.765 41.655 36.775 ;
        RECT 46.620 36.765 46.990 36.775 ;
        RECT 51.945 36.765 52.315 36.775 ;
        RECT 57.280 36.765 57.650 36.775 ;
        RECT 62.605 36.765 62.975 36.775 ;
        RECT 67.940 36.765 68.310 36.775 ;
        RECT 73.265 36.765 73.635 36.775 ;
        RECT 78.600 36.765 78.970 36.775 ;
        RECT 83.925 36.765 84.295 36.775 ;
        RECT 89.260 36.765 89.630 36.775 ;
        RECT 94.585 36.765 94.955 36.775 ;
        RECT 99.920 36.765 100.290 36.775 ;
        RECT 105.245 36.765 105.615 36.775 ;
        RECT 110.580 36.765 110.950 36.775 ;
        RECT 115.905 36.765 116.275 36.775 ;
        RECT 121.240 36.765 121.610 36.775 ;
        RECT 28.030 35.085 28.310 35.455 ;
        RECT 27.655 33.145 27.935 33.515 ;
        RECT 27.270 30.815 27.550 31.185 ;
        RECT 26.895 26.900 27.175 27.270 ;
        RECT 26.515 25.610 26.795 25.980 ;
        RECT 26.565 22.360 26.745 25.610 ;
        RECT 26.945 25.015 27.125 26.900 ;
        RECT 26.905 23.905 27.165 25.015 ;
        RECT 26.945 23.650 27.125 23.905 ;
        RECT 26.890 23.280 27.170 23.650 ;
        RECT 26.945 23.220 27.125 23.280 ;
        RECT 26.515 21.990 26.795 22.360 ;
        RECT 26.565 20.290 26.745 21.990 ;
        RECT 26.525 19.185 26.785 20.290 ;
        RECT 26.565 19.150 26.745 19.185 ;
        RECT 27.325 18.445 27.505 30.815 ;
        RECT 27.705 29.895 27.885 33.145 ;
        RECT 27.655 29.525 27.935 29.895 ;
        RECT 27.705 19.735 27.885 29.525 ;
        RECT 28.085 29.250 28.265 35.085 ;
        RECT 28.465 34.160 28.645 36.415 ;
        RECT 36.785 35.100 37.155 35.110 ;
        RECT 42.120 35.100 42.490 35.110 ;
        RECT 47.445 35.100 47.815 35.110 ;
        RECT 52.780 35.100 53.150 35.110 ;
        RECT 58.105 35.100 58.475 35.110 ;
        RECT 63.440 35.100 63.810 35.110 ;
        RECT 68.765 35.100 69.135 35.110 ;
        RECT 74.100 35.100 74.470 35.110 ;
        RECT 79.425 35.100 79.795 35.110 ;
        RECT 84.760 35.100 85.130 35.110 ;
        RECT 90.085 35.100 90.455 35.110 ;
        RECT 95.420 35.100 95.790 35.110 ;
        RECT 100.745 35.100 101.115 35.110 ;
        RECT 106.080 35.100 106.450 35.110 ;
        RECT 111.405 35.100 111.775 35.110 ;
        RECT 116.740 35.100 117.110 35.110 ;
        RECT 36.785 34.840 37.810 35.100 ;
        RECT 36.785 34.830 37.155 34.840 ;
        RECT 38.105 34.810 39.655 35.090 ;
        RECT 41.285 35.005 41.655 35.015 ;
        RECT 39.375 34.455 39.655 34.810 ;
        RECT 40.630 34.745 41.655 35.005 ;
        RECT 42.120 34.840 43.145 35.100 ;
        RECT 42.120 34.830 42.490 34.840 ;
        RECT 43.440 34.810 44.990 35.090 ;
        RECT 46.620 35.005 46.990 35.015 ;
        RECT 41.285 34.735 41.655 34.745 ;
        RECT 44.710 34.455 44.990 34.810 ;
        RECT 45.965 34.745 46.990 35.005 ;
        RECT 47.445 34.840 48.470 35.100 ;
        RECT 47.445 34.830 47.815 34.840 ;
        RECT 48.765 34.810 50.315 35.090 ;
        RECT 51.945 35.005 52.315 35.015 ;
        RECT 46.620 34.735 46.990 34.745 ;
        RECT 50.035 34.455 50.315 34.810 ;
        RECT 51.290 34.745 52.315 35.005 ;
        RECT 52.780 34.840 53.805 35.100 ;
        RECT 52.780 34.830 53.150 34.840 ;
        RECT 54.100 34.810 55.650 35.090 ;
        RECT 57.280 35.005 57.650 35.015 ;
        RECT 51.945 34.735 52.315 34.745 ;
        RECT 55.370 34.455 55.650 34.810 ;
        RECT 56.625 34.745 57.650 35.005 ;
        RECT 58.105 34.840 59.130 35.100 ;
        RECT 58.105 34.830 58.475 34.840 ;
        RECT 59.425 34.810 60.975 35.090 ;
        RECT 62.605 35.005 62.975 35.015 ;
        RECT 57.280 34.735 57.650 34.745 ;
        RECT 60.695 34.455 60.975 34.810 ;
        RECT 61.950 34.745 62.975 35.005 ;
        RECT 63.440 34.840 64.465 35.100 ;
        RECT 63.440 34.830 63.810 34.840 ;
        RECT 64.760 34.810 66.310 35.090 ;
        RECT 67.940 35.005 68.310 35.015 ;
        RECT 62.605 34.735 62.975 34.745 ;
        RECT 66.030 34.455 66.310 34.810 ;
        RECT 67.285 34.745 68.310 35.005 ;
        RECT 68.765 34.840 69.790 35.100 ;
        RECT 68.765 34.830 69.135 34.840 ;
        RECT 70.085 34.810 71.635 35.090 ;
        RECT 73.265 35.005 73.635 35.015 ;
        RECT 67.940 34.735 68.310 34.745 ;
        RECT 71.355 34.455 71.635 34.810 ;
        RECT 72.610 34.745 73.635 35.005 ;
        RECT 74.100 34.840 75.125 35.100 ;
        RECT 74.100 34.830 74.470 34.840 ;
        RECT 75.420 34.810 76.970 35.090 ;
        RECT 78.600 35.005 78.970 35.015 ;
        RECT 73.265 34.735 73.635 34.745 ;
        RECT 76.690 34.455 76.970 34.810 ;
        RECT 77.945 34.745 78.970 35.005 ;
        RECT 79.425 34.840 80.450 35.100 ;
        RECT 79.425 34.830 79.795 34.840 ;
        RECT 80.745 34.810 82.295 35.090 ;
        RECT 83.925 35.005 84.295 35.015 ;
        RECT 78.600 34.735 78.970 34.745 ;
        RECT 82.015 34.455 82.295 34.810 ;
        RECT 83.270 34.745 84.295 35.005 ;
        RECT 84.760 34.840 85.785 35.100 ;
        RECT 84.760 34.830 85.130 34.840 ;
        RECT 86.080 34.810 87.630 35.090 ;
        RECT 89.260 35.005 89.630 35.015 ;
        RECT 83.925 34.735 84.295 34.745 ;
        RECT 87.350 34.455 87.630 34.810 ;
        RECT 88.605 34.745 89.630 35.005 ;
        RECT 90.085 34.840 91.110 35.100 ;
        RECT 90.085 34.830 90.455 34.840 ;
        RECT 91.405 34.810 92.955 35.090 ;
        RECT 94.585 35.005 94.955 35.015 ;
        RECT 89.260 34.735 89.630 34.745 ;
        RECT 92.675 34.455 92.955 34.810 ;
        RECT 93.930 34.745 94.955 35.005 ;
        RECT 95.420 34.840 96.445 35.100 ;
        RECT 95.420 34.830 95.790 34.840 ;
        RECT 96.740 34.810 98.290 35.090 ;
        RECT 99.920 35.005 100.290 35.015 ;
        RECT 94.585 34.735 94.955 34.745 ;
        RECT 98.010 34.455 98.290 34.810 ;
        RECT 99.265 34.745 100.290 35.005 ;
        RECT 100.745 34.840 101.770 35.100 ;
        RECT 100.745 34.830 101.115 34.840 ;
        RECT 102.065 34.810 103.615 35.090 ;
        RECT 105.245 35.005 105.615 35.015 ;
        RECT 99.920 34.735 100.290 34.745 ;
        RECT 103.335 34.455 103.615 34.810 ;
        RECT 104.590 34.745 105.615 35.005 ;
        RECT 106.080 34.840 107.105 35.100 ;
        RECT 106.080 34.830 106.450 34.840 ;
        RECT 107.400 34.810 108.950 35.090 ;
        RECT 110.580 35.005 110.950 35.015 ;
        RECT 105.245 34.735 105.615 34.745 ;
        RECT 108.670 34.455 108.950 34.810 ;
        RECT 109.925 34.745 110.950 35.005 ;
        RECT 111.405 34.840 112.430 35.100 ;
        RECT 111.405 34.830 111.775 34.840 ;
        RECT 112.725 34.810 114.275 35.090 ;
        RECT 115.905 35.005 116.275 35.015 ;
        RECT 110.580 34.735 110.950 34.745 ;
        RECT 113.995 34.455 114.275 34.810 ;
        RECT 115.250 34.745 116.275 35.005 ;
        RECT 116.740 34.840 117.765 35.100 ;
        RECT 116.740 34.830 117.110 34.840 ;
        RECT 118.060 34.810 119.610 35.090 ;
        RECT 121.240 35.005 121.610 35.015 ;
        RECT 115.905 34.735 116.275 34.745 ;
        RECT 119.330 34.455 119.610 34.810 ;
        RECT 120.585 34.745 121.610 35.005 ;
        RECT 121.240 34.735 121.610 34.745 ;
        RECT 34.005 34.450 34.400 34.455 ;
        RECT 33.390 34.170 35.160 34.450 ;
        RECT 38.715 34.170 39.110 34.450 ;
        RECT 39.330 34.175 39.725 34.455 ;
        RECT 40.015 34.170 40.485 34.450 ;
        RECT 44.050 34.170 44.445 34.450 ;
        RECT 44.665 34.175 45.060 34.455 ;
        RECT 45.350 34.170 45.820 34.450 ;
        RECT 49.375 34.170 49.770 34.450 ;
        RECT 49.990 34.175 50.385 34.455 ;
        RECT 50.675 34.170 51.145 34.450 ;
        RECT 54.710 34.170 55.105 34.450 ;
        RECT 55.325 34.175 55.720 34.455 ;
        RECT 56.010 34.170 56.480 34.450 ;
        RECT 60.035 34.170 60.430 34.450 ;
        RECT 60.650 34.175 61.045 34.455 ;
        RECT 61.335 34.170 61.805 34.450 ;
        RECT 65.370 34.170 65.765 34.450 ;
        RECT 65.985 34.175 66.380 34.455 ;
        RECT 66.670 34.170 67.140 34.450 ;
        RECT 70.695 34.170 71.090 34.450 ;
        RECT 71.310 34.175 71.705 34.455 ;
        RECT 71.995 34.170 72.465 34.450 ;
        RECT 76.030 34.170 76.425 34.450 ;
        RECT 76.645 34.175 77.040 34.455 ;
        RECT 77.330 34.170 77.800 34.450 ;
        RECT 81.355 34.170 81.750 34.450 ;
        RECT 81.970 34.175 82.365 34.455 ;
        RECT 82.655 34.170 83.125 34.450 ;
        RECT 86.690 34.170 87.085 34.450 ;
        RECT 87.305 34.175 87.700 34.455 ;
        RECT 87.990 34.170 88.460 34.450 ;
        RECT 92.015 34.170 92.410 34.450 ;
        RECT 92.630 34.175 93.025 34.455 ;
        RECT 93.315 34.170 93.785 34.450 ;
        RECT 97.350 34.170 97.745 34.450 ;
        RECT 97.965 34.175 98.360 34.455 ;
        RECT 98.650 34.170 99.120 34.450 ;
        RECT 102.675 34.170 103.070 34.450 ;
        RECT 103.290 34.175 103.685 34.455 ;
        RECT 103.975 34.170 104.445 34.450 ;
        RECT 108.010 34.170 108.405 34.450 ;
        RECT 108.625 34.175 109.020 34.455 ;
        RECT 109.310 34.170 109.780 34.450 ;
        RECT 113.335 34.170 113.730 34.450 ;
        RECT 113.950 34.175 114.345 34.455 ;
        RECT 114.635 34.170 115.105 34.450 ;
        RECT 118.670 34.170 119.065 34.450 ;
        RECT 119.285 34.175 119.680 34.455 ;
        RECT 124.610 34.450 125.005 34.455 ;
        RECT 119.970 34.170 120.440 34.450 ;
        RECT 123.995 34.170 125.765 34.450 ;
        RECT 28.415 33.790 28.695 34.160 ;
        RECT 36.785 33.800 37.155 33.810 ;
        RECT 42.120 33.800 42.490 33.810 ;
        RECT 47.445 33.800 47.815 33.810 ;
        RECT 52.780 33.800 53.150 33.810 ;
        RECT 58.105 33.800 58.475 33.810 ;
        RECT 63.440 33.800 63.810 33.810 ;
        RECT 68.765 33.800 69.135 33.810 ;
        RECT 74.100 33.800 74.470 33.810 ;
        RECT 79.425 33.800 79.795 33.810 ;
        RECT 84.760 33.800 85.130 33.810 ;
        RECT 90.085 33.800 90.455 33.810 ;
        RECT 95.420 33.800 95.790 33.810 ;
        RECT 100.745 33.800 101.115 33.810 ;
        RECT 106.080 33.800 106.450 33.810 ;
        RECT 111.405 33.800 111.775 33.810 ;
        RECT 116.740 33.800 117.110 33.810 ;
        RECT 28.465 30.540 28.645 33.790 ;
        RECT 36.785 33.540 37.860 33.800 ;
        RECT 42.120 33.540 43.195 33.800 ;
        RECT 47.445 33.540 48.520 33.800 ;
        RECT 52.780 33.540 53.855 33.800 ;
        RECT 58.105 33.540 59.180 33.800 ;
        RECT 63.440 33.540 64.515 33.800 ;
        RECT 68.765 33.540 69.840 33.800 ;
        RECT 74.100 33.540 75.175 33.800 ;
        RECT 79.425 33.540 80.500 33.800 ;
        RECT 84.760 33.540 85.835 33.800 ;
        RECT 90.085 33.540 91.160 33.800 ;
        RECT 95.420 33.540 96.495 33.800 ;
        RECT 100.745 33.540 101.820 33.800 ;
        RECT 106.080 33.540 107.155 33.800 ;
        RECT 111.405 33.540 112.480 33.800 ;
        RECT 116.740 33.540 117.815 33.800 ;
        RECT 36.785 33.530 37.155 33.540 ;
        RECT 42.120 33.530 42.490 33.540 ;
        RECT 47.445 33.530 47.815 33.540 ;
        RECT 52.780 33.530 53.150 33.540 ;
        RECT 58.105 33.530 58.475 33.540 ;
        RECT 63.440 33.530 63.810 33.540 ;
        RECT 68.765 33.530 69.135 33.540 ;
        RECT 74.100 33.530 74.470 33.540 ;
        RECT 79.425 33.530 79.795 33.540 ;
        RECT 84.760 33.530 85.130 33.540 ;
        RECT 90.085 33.530 90.455 33.540 ;
        RECT 95.420 33.530 95.790 33.540 ;
        RECT 100.745 33.530 101.115 33.540 ;
        RECT 106.080 33.530 106.450 33.540 ;
        RECT 111.405 33.530 111.775 33.540 ;
        RECT 116.740 33.530 117.110 33.540 ;
        RECT 41.290 33.170 41.660 33.180 ;
        RECT 46.625 33.170 46.995 33.180 ;
        RECT 51.950 33.170 52.320 33.180 ;
        RECT 57.285 33.170 57.655 33.180 ;
        RECT 62.610 33.170 62.980 33.180 ;
        RECT 67.945 33.170 68.315 33.180 ;
        RECT 73.270 33.170 73.640 33.180 ;
        RECT 78.605 33.170 78.975 33.180 ;
        RECT 83.930 33.170 84.300 33.180 ;
        RECT 89.265 33.170 89.635 33.180 ;
        RECT 94.590 33.170 94.960 33.180 ;
        RECT 99.925 33.170 100.295 33.180 ;
        RECT 105.250 33.170 105.620 33.180 ;
        RECT 110.585 33.170 110.955 33.180 ;
        RECT 115.910 33.170 116.280 33.180 ;
        RECT 121.245 33.170 121.615 33.180 ;
        RECT 40.630 32.910 41.660 33.170 ;
        RECT 45.965 32.910 46.995 33.170 ;
        RECT 51.290 32.910 52.320 33.170 ;
        RECT 56.625 32.910 57.655 33.170 ;
        RECT 61.950 32.910 62.980 33.170 ;
        RECT 67.285 32.910 68.315 33.170 ;
        RECT 72.610 32.910 73.640 33.170 ;
        RECT 77.945 32.910 78.975 33.170 ;
        RECT 83.270 32.910 84.300 33.170 ;
        RECT 88.605 32.910 89.635 33.170 ;
        RECT 93.930 32.910 94.960 33.170 ;
        RECT 99.265 32.910 100.295 33.170 ;
        RECT 104.590 32.910 105.620 33.170 ;
        RECT 109.925 32.910 110.955 33.170 ;
        RECT 115.250 32.910 116.280 33.170 ;
        RECT 120.585 32.910 121.615 33.170 ;
        RECT 41.290 32.900 41.660 32.910 ;
        RECT 46.625 32.900 46.995 32.910 ;
        RECT 51.950 32.900 52.320 32.910 ;
        RECT 57.285 32.900 57.655 32.910 ;
        RECT 62.610 32.900 62.980 32.910 ;
        RECT 67.945 32.900 68.315 32.910 ;
        RECT 73.270 32.900 73.640 32.910 ;
        RECT 78.605 32.900 78.975 32.910 ;
        RECT 83.930 32.900 84.300 32.910 ;
        RECT 89.265 32.900 89.635 32.910 ;
        RECT 94.590 32.900 94.960 32.910 ;
        RECT 99.925 32.900 100.295 32.910 ;
        RECT 105.250 32.900 105.620 32.910 ;
        RECT 110.585 32.900 110.955 32.910 ;
        RECT 115.910 32.900 116.280 32.910 ;
        RECT 121.245 32.900 121.615 32.910 ;
        RECT 36.790 31.435 37.160 31.445 ;
        RECT 42.125 31.435 42.495 31.445 ;
        RECT 47.450 31.435 47.820 31.445 ;
        RECT 52.785 31.435 53.155 31.445 ;
        RECT 58.110 31.435 58.480 31.445 ;
        RECT 63.445 31.435 63.815 31.445 ;
        RECT 68.770 31.435 69.140 31.445 ;
        RECT 74.105 31.435 74.475 31.445 ;
        RECT 79.430 31.435 79.800 31.445 ;
        RECT 84.765 31.435 85.135 31.445 ;
        RECT 90.090 31.435 90.460 31.445 ;
        RECT 95.425 31.435 95.795 31.445 ;
        RECT 100.750 31.435 101.120 31.445 ;
        RECT 106.085 31.435 106.455 31.445 ;
        RECT 111.410 31.435 111.780 31.445 ;
        RECT 116.745 31.435 117.115 31.445 ;
        RECT 36.790 31.175 37.810 31.435 ;
        RECT 42.125 31.175 43.145 31.435 ;
        RECT 47.450 31.175 48.470 31.435 ;
        RECT 52.785 31.175 53.805 31.435 ;
        RECT 58.110 31.175 59.130 31.435 ;
        RECT 63.445 31.175 64.465 31.435 ;
        RECT 68.770 31.175 69.790 31.435 ;
        RECT 74.105 31.175 75.125 31.435 ;
        RECT 79.430 31.175 80.450 31.435 ;
        RECT 84.765 31.175 85.785 31.435 ;
        RECT 90.090 31.175 91.110 31.435 ;
        RECT 95.425 31.175 96.445 31.435 ;
        RECT 100.750 31.175 101.770 31.435 ;
        RECT 106.085 31.175 107.105 31.435 ;
        RECT 111.410 31.175 112.430 31.435 ;
        RECT 116.745 31.175 117.765 31.435 ;
        RECT 36.790 31.165 37.160 31.175 ;
        RECT 42.125 31.165 42.495 31.175 ;
        RECT 47.450 31.165 47.820 31.175 ;
        RECT 52.785 31.165 53.155 31.175 ;
        RECT 58.110 31.165 58.480 31.175 ;
        RECT 63.445 31.165 63.815 31.175 ;
        RECT 68.770 31.165 69.140 31.175 ;
        RECT 74.105 31.165 74.475 31.175 ;
        RECT 79.430 31.165 79.800 31.175 ;
        RECT 84.765 31.165 85.135 31.175 ;
        RECT 90.090 31.165 90.460 31.175 ;
        RECT 95.425 31.165 95.795 31.175 ;
        RECT 100.750 31.165 101.120 31.175 ;
        RECT 106.085 31.165 106.455 31.175 ;
        RECT 111.410 31.165 111.780 31.175 ;
        RECT 116.745 31.165 117.115 31.175 ;
        RECT 28.415 30.170 28.695 30.540 ;
        RECT 38.105 30.520 39.655 30.800 ;
        RECT 41.285 30.785 41.655 30.795 ;
        RECT 40.580 30.525 41.655 30.785 ;
        RECT 28.035 28.880 28.315 29.250 ;
        RECT 28.085 26.625 28.265 28.880 ;
        RECT 28.465 27.920 28.645 30.170 ;
        RECT 39.375 30.090 39.655 30.520 ;
        RECT 41.285 30.515 41.655 30.525 ;
        RECT 43.440 30.520 44.990 30.800 ;
        RECT 46.620 30.785 46.990 30.795 ;
        RECT 45.915 30.525 46.990 30.785 ;
        RECT 44.710 30.090 44.990 30.520 ;
        RECT 46.620 30.515 46.990 30.525 ;
        RECT 48.765 30.520 50.315 30.800 ;
        RECT 51.945 30.785 52.315 30.795 ;
        RECT 51.240 30.525 52.315 30.785 ;
        RECT 50.035 30.090 50.315 30.520 ;
        RECT 51.945 30.515 52.315 30.525 ;
        RECT 54.100 30.520 55.650 30.800 ;
        RECT 57.280 30.785 57.650 30.795 ;
        RECT 56.575 30.525 57.650 30.785 ;
        RECT 55.370 30.090 55.650 30.520 ;
        RECT 57.280 30.515 57.650 30.525 ;
        RECT 59.425 30.520 60.975 30.800 ;
        RECT 62.605 30.785 62.975 30.795 ;
        RECT 61.900 30.525 62.975 30.785 ;
        RECT 60.695 30.090 60.975 30.520 ;
        RECT 62.605 30.515 62.975 30.525 ;
        RECT 64.760 30.520 66.310 30.800 ;
        RECT 67.940 30.785 68.310 30.795 ;
        RECT 67.235 30.525 68.310 30.785 ;
        RECT 66.030 30.090 66.310 30.520 ;
        RECT 67.940 30.515 68.310 30.525 ;
        RECT 70.085 30.520 71.635 30.800 ;
        RECT 73.265 30.785 73.635 30.795 ;
        RECT 72.560 30.525 73.635 30.785 ;
        RECT 71.355 30.090 71.635 30.520 ;
        RECT 73.265 30.515 73.635 30.525 ;
        RECT 75.420 30.520 76.970 30.800 ;
        RECT 78.600 30.785 78.970 30.795 ;
        RECT 77.895 30.525 78.970 30.785 ;
        RECT 76.690 30.090 76.970 30.520 ;
        RECT 78.600 30.515 78.970 30.525 ;
        RECT 80.745 30.520 82.295 30.800 ;
        RECT 83.925 30.785 84.295 30.795 ;
        RECT 83.220 30.525 84.295 30.785 ;
        RECT 82.015 30.090 82.295 30.520 ;
        RECT 83.925 30.515 84.295 30.525 ;
        RECT 86.080 30.520 87.630 30.800 ;
        RECT 89.260 30.785 89.630 30.795 ;
        RECT 88.555 30.525 89.630 30.785 ;
        RECT 87.350 30.090 87.630 30.520 ;
        RECT 89.260 30.515 89.630 30.525 ;
        RECT 91.405 30.520 92.955 30.800 ;
        RECT 94.585 30.785 94.955 30.795 ;
        RECT 93.880 30.525 94.955 30.785 ;
        RECT 92.675 30.090 92.955 30.520 ;
        RECT 94.585 30.515 94.955 30.525 ;
        RECT 96.740 30.520 98.290 30.800 ;
        RECT 99.920 30.785 100.290 30.795 ;
        RECT 99.215 30.525 100.290 30.785 ;
        RECT 98.010 30.090 98.290 30.520 ;
        RECT 99.920 30.515 100.290 30.525 ;
        RECT 102.065 30.520 103.615 30.800 ;
        RECT 105.245 30.785 105.615 30.795 ;
        RECT 104.540 30.525 105.615 30.785 ;
        RECT 103.335 30.090 103.615 30.520 ;
        RECT 105.245 30.515 105.615 30.525 ;
        RECT 107.400 30.520 108.950 30.800 ;
        RECT 110.580 30.785 110.950 30.795 ;
        RECT 109.875 30.525 110.950 30.785 ;
        RECT 108.670 30.090 108.950 30.520 ;
        RECT 110.580 30.515 110.950 30.525 ;
        RECT 112.725 30.520 114.275 30.800 ;
        RECT 115.905 30.785 116.275 30.795 ;
        RECT 115.200 30.525 116.275 30.785 ;
        RECT 113.995 30.090 114.275 30.520 ;
        RECT 115.905 30.515 116.275 30.525 ;
        RECT 118.060 30.520 119.610 30.800 ;
        RECT 121.240 30.785 121.610 30.795 ;
        RECT 120.535 30.525 121.610 30.785 ;
        RECT 119.330 30.090 119.610 30.520 ;
        RECT 121.240 30.515 121.610 30.525 ;
        RECT 32.625 29.810 34.390 30.090 ;
        RECT 37.950 29.810 38.470 30.090 ;
        RECT 38.715 29.810 39.110 30.090 ;
        RECT 39.330 29.810 39.715 30.090 ;
        RECT 43.285 29.810 43.805 30.090 ;
        RECT 44.050 29.810 44.445 30.090 ;
        RECT 44.665 29.810 45.050 30.090 ;
        RECT 48.610 29.810 49.130 30.090 ;
        RECT 49.375 29.810 49.770 30.090 ;
        RECT 49.990 29.810 50.375 30.090 ;
        RECT 53.945 29.810 54.465 30.090 ;
        RECT 54.710 29.810 55.105 30.090 ;
        RECT 55.325 29.810 55.710 30.090 ;
        RECT 59.270 29.810 59.790 30.090 ;
        RECT 60.035 29.810 60.430 30.090 ;
        RECT 60.650 29.810 61.035 30.090 ;
        RECT 64.605 29.810 65.125 30.090 ;
        RECT 65.370 29.810 65.765 30.090 ;
        RECT 65.985 29.810 66.370 30.090 ;
        RECT 69.930 29.810 70.450 30.090 ;
        RECT 70.695 29.810 71.090 30.090 ;
        RECT 71.310 29.810 71.695 30.090 ;
        RECT 75.265 29.810 75.785 30.090 ;
        RECT 76.030 29.810 76.425 30.090 ;
        RECT 76.645 29.810 77.030 30.090 ;
        RECT 80.590 29.810 81.110 30.090 ;
        RECT 81.355 29.810 81.750 30.090 ;
        RECT 81.970 29.810 82.355 30.090 ;
        RECT 85.925 29.810 86.445 30.090 ;
        RECT 86.690 29.810 87.085 30.090 ;
        RECT 87.305 29.810 87.690 30.090 ;
        RECT 91.250 29.810 91.770 30.090 ;
        RECT 92.015 29.810 92.410 30.090 ;
        RECT 92.630 29.810 93.015 30.090 ;
        RECT 96.585 29.810 97.105 30.090 ;
        RECT 97.350 29.810 97.745 30.090 ;
        RECT 97.965 29.810 98.350 30.090 ;
        RECT 101.910 29.810 102.430 30.090 ;
        RECT 102.675 29.810 103.070 30.090 ;
        RECT 103.290 29.810 103.675 30.090 ;
        RECT 107.245 29.810 107.765 30.090 ;
        RECT 108.010 29.810 108.405 30.090 ;
        RECT 108.625 29.810 109.010 30.090 ;
        RECT 112.570 29.810 113.090 30.090 ;
        RECT 113.335 29.810 113.730 30.090 ;
        RECT 113.950 29.810 114.335 30.090 ;
        RECT 117.905 29.810 118.425 30.090 ;
        RECT 118.670 29.810 119.065 30.090 ;
        RECT 119.285 29.810 119.670 30.090 ;
        RECT 123.230 29.810 124.995 30.090 ;
        RECT 36.785 29.590 37.155 29.600 ;
        RECT 42.120 29.590 42.490 29.600 ;
        RECT 47.445 29.590 47.815 29.600 ;
        RECT 52.780 29.590 53.150 29.600 ;
        RECT 58.105 29.590 58.475 29.600 ;
        RECT 63.440 29.590 63.810 29.600 ;
        RECT 68.765 29.590 69.135 29.600 ;
        RECT 74.100 29.590 74.470 29.600 ;
        RECT 79.425 29.590 79.795 29.600 ;
        RECT 84.760 29.590 85.130 29.600 ;
        RECT 90.085 29.590 90.455 29.600 ;
        RECT 95.420 29.590 95.790 29.600 ;
        RECT 100.745 29.590 101.115 29.600 ;
        RECT 106.080 29.590 106.450 29.600 ;
        RECT 111.405 29.590 111.775 29.600 ;
        RECT 116.740 29.590 117.110 29.600 ;
        RECT 36.785 29.330 37.810 29.590 ;
        RECT 41.285 29.500 41.655 29.510 ;
        RECT 36.785 29.320 37.155 29.330 ;
        RECT 40.630 29.240 41.655 29.500 ;
        RECT 42.120 29.330 43.145 29.590 ;
        RECT 46.620 29.500 46.990 29.510 ;
        RECT 42.120 29.320 42.490 29.330 ;
        RECT 45.965 29.240 46.990 29.500 ;
        RECT 47.445 29.330 48.470 29.590 ;
        RECT 51.945 29.500 52.315 29.510 ;
        RECT 47.445 29.320 47.815 29.330 ;
        RECT 51.290 29.240 52.315 29.500 ;
        RECT 52.780 29.330 53.805 29.590 ;
        RECT 57.280 29.500 57.650 29.510 ;
        RECT 52.780 29.320 53.150 29.330 ;
        RECT 56.625 29.240 57.650 29.500 ;
        RECT 58.105 29.330 59.130 29.590 ;
        RECT 62.605 29.500 62.975 29.510 ;
        RECT 58.105 29.320 58.475 29.330 ;
        RECT 61.950 29.240 62.975 29.500 ;
        RECT 63.440 29.330 64.465 29.590 ;
        RECT 67.940 29.500 68.310 29.510 ;
        RECT 63.440 29.320 63.810 29.330 ;
        RECT 67.285 29.240 68.310 29.500 ;
        RECT 68.765 29.330 69.790 29.590 ;
        RECT 73.265 29.500 73.635 29.510 ;
        RECT 68.765 29.320 69.135 29.330 ;
        RECT 72.610 29.240 73.635 29.500 ;
        RECT 74.100 29.330 75.125 29.590 ;
        RECT 78.600 29.500 78.970 29.510 ;
        RECT 74.100 29.320 74.470 29.330 ;
        RECT 77.945 29.240 78.970 29.500 ;
        RECT 79.425 29.330 80.450 29.590 ;
        RECT 83.925 29.500 84.295 29.510 ;
        RECT 79.425 29.320 79.795 29.330 ;
        RECT 83.270 29.240 84.295 29.500 ;
        RECT 84.760 29.330 85.785 29.590 ;
        RECT 89.260 29.500 89.630 29.510 ;
        RECT 84.760 29.320 85.130 29.330 ;
        RECT 88.605 29.240 89.630 29.500 ;
        RECT 90.085 29.330 91.110 29.590 ;
        RECT 94.585 29.500 94.955 29.510 ;
        RECT 90.085 29.320 90.455 29.330 ;
        RECT 93.930 29.240 94.955 29.500 ;
        RECT 95.420 29.330 96.445 29.590 ;
        RECT 99.920 29.500 100.290 29.510 ;
        RECT 95.420 29.320 95.790 29.330 ;
        RECT 99.265 29.240 100.290 29.500 ;
        RECT 100.745 29.330 101.770 29.590 ;
        RECT 105.245 29.500 105.615 29.510 ;
        RECT 100.745 29.320 101.115 29.330 ;
        RECT 104.590 29.240 105.615 29.500 ;
        RECT 106.080 29.330 107.105 29.590 ;
        RECT 110.580 29.500 110.950 29.510 ;
        RECT 106.080 29.320 106.450 29.330 ;
        RECT 109.925 29.240 110.950 29.500 ;
        RECT 111.405 29.330 112.430 29.590 ;
        RECT 115.905 29.500 116.275 29.510 ;
        RECT 111.405 29.320 111.775 29.330 ;
        RECT 115.250 29.240 116.275 29.500 ;
        RECT 116.740 29.330 117.765 29.590 ;
        RECT 121.240 29.500 121.610 29.510 ;
        RECT 116.740 29.320 117.110 29.330 ;
        RECT 120.585 29.240 121.610 29.500 ;
        RECT 41.285 29.230 41.655 29.240 ;
        RECT 46.620 29.230 46.990 29.240 ;
        RECT 51.945 29.230 52.315 29.240 ;
        RECT 57.280 29.230 57.650 29.240 ;
        RECT 62.605 29.230 62.975 29.240 ;
        RECT 67.940 29.230 68.310 29.240 ;
        RECT 73.265 29.230 73.635 29.240 ;
        RECT 78.600 29.230 78.970 29.240 ;
        RECT 83.925 29.230 84.295 29.240 ;
        RECT 89.260 29.230 89.630 29.240 ;
        RECT 94.585 29.230 94.955 29.240 ;
        RECT 99.920 29.230 100.290 29.240 ;
        RECT 105.245 29.230 105.615 29.240 ;
        RECT 110.580 29.230 110.950 29.240 ;
        RECT 115.905 29.230 116.275 29.240 ;
        RECT 121.240 29.230 121.610 29.240 ;
        RECT 28.410 27.550 28.690 27.920 ;
        RECT 36.785 27.565 37.155 27.575 ;
        RECT 42.120 27.565 42.490 27.575 ;
        RECT 47.445 27.565 47.815 27.575 ;
        RECT 52.780 27.565 53.150 27.575 ;
        RECT 58.105 27.565 58.475 27.575 ;
        RECT 63.440 27.565 63.810 27.575 ;
        RECT 68.765 27.565 69.135 27.575 ;
        RECT 74.100 27.565 74.470 27.575 ;
        RECT 79.425 27.565 79.795 27.575 ;
        RECT 84.760 27.565 85.130 27.575 ;
        RECT 90.085 27.565 90.455 27.575 ;
        RECT 95.420 27.565 95.790 27.575 ;
        RECT 100.745 27.565 101.115 27.575 ;
        RECT 106.080 27.565 106.450 27.575 ;
        RECT 111.405 27.565 111.775 27.575 ;
        RECT 116.740 27.565 117.110 27.575 ;
        RECT 28.035 26.255 28.315 26.625 ;
        RECT 28.085 23.005 28.265 26.255 ;
        RECT 28.035 22.635 28.315 23.005 ;
        RECT 28.085 20.385 28.265 22.635 ;
        RECT 28.465 21.715 28.645 27.550 ;
        RECT 36.785 27.305 37.810 27.565 ;
        RECT 41.285 27.470 41.655 27.480 ;
        RECT 36.785 27.295 37.155 27.305 ;
        RECT 40.630 27.210 41.655 27.470 ;
        RECT 42.120 27.305 43.145 27.565 ;
        RECT 46.620 27.470 46.990 27.480 ;
        RECT 42.120 27.295 42.490 27.305 ;
        RECT 45.965 27.210 46.990 27.470 ;
        RECT 47.445 27.305 48.470 27.565 ;
        RECT 51.945 27.470 52.315 27.480 ;
        RECT 47.445 27.295 47.815 27.305 ;
        RECT 51.290 27.210 52.315 27.470 ;
        RECT 52.780 27.305 53.805 27.565 ;
        RECT 57.280 27.470 57.650 27.480 ;
        RECT 52.780 27.295 53.150 27.305 ;
        RECT 56.625 27.210 57.650 27.470 ;
        RECT 58.105 27.305 59.130 27.565 ;
        RECT 62.605 27.470 62.975 27.480 ;
        RECT 58.105 27.295 58.475 27.305 ;
        RECT 61.950 27.210 62.975 27.470 ;
        RECT 63.440 27.305 64.465 27.565 ;
        RECT 67.940 27.470 68.310 27.480 ;
        RECT 63.440 27.295 63.810 27.305 ;
        RECT 67.285 27.210 68.310 27.470 ;
        RECT 68.765 27.305 69.790 27.565 ;
        RECT 73.265 27.470 73.635 27.480 ;
        RECT 68.765 27.295 69.135 27.305 ;
        RECT 72.610 27.210 73.635 27.470 ;
        RECT 74.100 27.305 75.125 27.565 ;
        RECT 78.600 27.470 78.970 27.480 ;
        RECT 74.100 27.295 74.470 27.305 ;
        RECT 77.945 27.210 78.970 27.470 ;
        RECT 79.425 27.305 80.450 27.565 ;
        RECT 83.925 27.470 84.295 27.480 ;
        RECT 79.425 27.295 79.795 27.305 ;
        RECT 83.270 27.210 84.295 27.470 ;
        RECT 84.760 27.305 85.785 27.565 ;
        RECT 89.260 27.470 89.630 27.480 ;
        RECT 84.760 27.295 85.130 27.305 ;
        RECT 88.605 27.210 89.630 27.470 ;
        RECT 90.085 27.305 91.110 27.565 ;
        RECT 94.585 27.470 94.955 27.480 ;
        RECT 90.085 27.295 90.455 27.305 ;
        RECT 93.930 27.210 94.955 27.470 ;
        RECT 95.420 27.305 96.445 27.565 ;
        RECT 99.920 27.470 100.290 27.480 ;
        RECT 95.420 27.295 95.790 27.305 ;
        RECT 99.265 27.210 100.290 27.470 ;
        RECT 100.745 27.305 101.770 27.565 ;
        RECT 105.245 27.470 105.615 27.480 ;
        RECT 100.745 27.295 101.115 27.305 ;
        RECT 104.590 27.210 105.615 27.470 ;
        RECT 106.080 27.305 107.105 27.565 ;
        RECT 110.580 27.470 110.950 27.480 ;
        RECT 106.080 27.295 106.450 27.305 ;
        RECT 109.925 27.210 110.950 27.470 ;
        RECT 111.405 27.305 112.430 27.565 ;
        RECT 115.905 27.470 116.275 27.480 ;
        RECT 111.405 27.295 111.775 27.305 ;
        RECT 115.250 27.210 116.275 27.470 ;
        RECT 116.740 27.305 117.765 27.565 ;
        RECT 121.240 27.470 121.610 27.480 ;
        RECT 116.740 27.295 117.110 27.305 ;
        RECT 120.585 27.210 121.610 27.470 ;
        RECT 41.285 27.200 41.655 27.210 ;
        RECT 46.620 27.200 46.990 27.210 ;
        RECT 51.945 27.200 52.315 27.210 ;
        RECT 57.280 27.200 57.650 27.210 ;
        RECT 62.605 27.200 62.975 27.210 ;
        RECT 67.940 27.200 68.310 27.210 ;
        RECT 73.265 27.200 73.635 27.210 ;
        RECT 78.600 27.200 78.970 27.210 ;
        RECT 83.925 27.200 84.295 27.210 ;
        RECT 89.260 27.200 89.630 27.210 ;
        RECT 94.585 27.200 94.955 27.210 ;
        RECT 99.920 27.200 100.290 27.210 ;
        RECT 105.245 27.200 105.615 27.210 ;
        RECT 110.580 27.200 110.950 27.210 ;
        RECT 115.905 27.200 116.275 27.210 ;
        RECT 121.240 27.200 121.610 27.210 ;
        RECT 34.005 26.915 34.400 26.920 ;
        RECT 33.390 26.635 35.160 26.915 ;
        RECT 38.715 26.635 39.110 26.915 ;
        RECT 39.330 26.640 39.725 26.920 ;
        RECT 39.385 26.330 39.645 26.640 ;
        RECT 40.030 26.635 40.485 26.915 ;
        RECT 44.050 26.635 44.445 26.915 ;
        RECT 44.665 26.640 45.060 26.920 ;
        RECT 44.720 26.330 44.980 26.640 ;
        RECT 45.365 26.635 45.820 26.915 ;
        RECT 49.375 26.635 49.770 26.915 ;
        RECT 49.990 26.640 50.385 26.920 ;
        RECT 50.045 26.330 50.305 26.640 ;
        RECT 50.690 26.635 51.145 26.915 ;
        RECT 54.710 26.635 55.105 26.915 ;
        RECT 55.325 26.640 55.720 26.920 ;
        RECT 55.380 26.330 55.640 26.640 ;
        RECT 56.025 26.635 56.480 26.915 ;
        RECT 60.035 26.635 60.430 26.915 ;
        RECT 60.650 26.640 61.045 26.920 ;
        RECT 60.705 26.330 60.965 26.640 ;
        RECT 61.350 26.635 61.805 26.915 ;
        RECT 65.370 26.635 65.765 26.915 ;
        RECT 65.985 26.640 66.380 26.920 ;
        RECT 66.040 26.330 66.300 26.640 ;
        RECT 66.685 26.635 67.140 26.915 ;
        RECT 70.695 26.635 71.090 26.915 ;
        RECT 71.310 26.640 71.705 26.920 ;
        RECT 71.365 26.330 71.625 26.640 ;
        RECT 72.010 26.635 72.465 26.915 ;
        RECT 76.030 26.635 76.425 26.915 ;
        RECT 76.645 26.640 77.040 26.920 ;
        RECT 76.700 26.330 76.960 26.640 ;
        RECT 77.345 26.635 77.800 26.915 ;
        RECT 81.355 26.635 81.750 26.915 ;
        RECT 81.970 26.640 82.365 26.920 ;
        RECT 82.025 26.330 82.285 26.640 ;
        RECT 82.670 26.635 83.125 26.915 ;
        RECT 86.690 26.635 87.085 26.915 ;
        RECT 87.305 26.640 87.700 26.920 ;
        RECT 87.360 26.330 87.620 26.640 ;
        RECT 88.005 26.635 88.460 26.915 ;
        RECT 92.015 26.635 92.410 26.915 ;
        RECT 92.630 26.640 93.025 26.920 ;
        RECT 92.685 26.330 92.945 26.640 ;
        RECT 93.330 26.635 93.785 26.915 ;
        RECT 97.350 26.635 97.745 26.915 ;
        RECT 97.965 26.640 98.360 26.920 ;
        RECT 98.020 26.330 98.280 26.640 ;
        RECT 98.665 26.635 99.120 26.915 ;
        RECT 102.675 26.635 103.070 26.915 ;
        RECT 103.290 26.640 103.685 26.920 ;
        RECT 103.345 26.330 103.605 26.640 ;
        RECT 103.990 26.635 104.445 26.915 ;
        RECT 108.010 26.635 108.405 26.915 ;
        RECT 108.625 26.640 109.020 26.920 ;
        RECT 108.680 26.330 108.940 26.640 ;
        RECT 109.325 26.635 109.780 26.915 ;
        RECT 113.335 26.635 113.730 26.915 ;
        RECT 113.950 26.640 114.345 26.920 ;
        RECT 114.005 26.330 114.265 26.640 ;
        RECT 114.650 26.635 115.105 26.915 ;
        RECT 118.670 26.635 119.065 26.915 ;
        RECT 119.285 26.640 119.680 26.920 ;
        RECT 124.610 26.915 125.005 26.920 ;
        RECT 119.340 26.330 119.600 26.640 ;
        RECT 119.985 26.635 120.440 26.915 ;
        RECT 123.995 26.635 125.765 26.915 ;
        RECT 36.785 26.265 37.155 26.275 ;
        RECT 36.785 26.005 37.860 26.265 ;
        RECT 39.385 26.050 41.015 26.330 ;
        RECT 42.120 26.265 42.490 26.275 ;
        RECT 42.120 26.005 43.195 26.265 ;
        RECT 44.720 26.050 46.350 26.330 ;
        RECT 47.445 26.265 47.815 26.275 ;
        RECT 47.445 26.005 48.520 26.265 ;
        RECT 50.045 26.050 51.675 26.330 ;
        RECT 52.780 26.265 53.150 26.275 ;
        RECT 52.780 26.005 53.855 26.265 ;
        RECT 55.380 26.050 57.010 26.330 ;
        RECT 58.105 26.265 58.475 26.275 ;
        RECT 58.105 26.005 59.180 26.265 ;
        RECT 60.705 26.050 62.335 26.330 ;
        RECT 63.440 26.265 63.810 26.275 ;
        RECT 63.440 26.005 64.515 26.265 ;
        RECT 66.040 26.050 67.670 26.330 ;
        RECT 68.765 26.265 69.135 26.275 ;
        RECT 68.765 26.005 69.840 26.265 ;
        RECT 71.365 26.050 72.995 26.330 ;
        RECT 74.100 26.265 74.470 26.275 ;
        RECT 74.100 26.005 75.175 26.265 ;
        RECT 76.700 26.050 78.330 26.330 ;
        RECT 79.425 26.265 79.795 26.275 ;
        RECT 79.425 26.005 80.500 26.265 ;
        RECT 82.025 26.050 83.655 26.330 ;
        RECT 84.760 26.265 85.130 26.275 ;
        RECT 84.760 26.005 85.835 26.265 ;
        RECT 87.360 26.050 88.990 26.330 ;
        RECT 90.085 26.265 90.455 26.275 ;
        RECT 90.085 26.005 91.160 26.265 ;
        RECT 92.685 26.050 94.315 26.330 ;
        RECT 95.420 26.265 95.790 26.275 ;
        RECT 95.420 26.005 96.495 26.265 ;
        RECT 98.020 26.050 99.650 26.330 ;
        RECT 100.745 26.265 101.115 26.275 ;
        RECT 100.745 26.005 101.820 26.265 ;
        RECT 103.345 26.050 104.975 26.330 ;
        RECT 106.080 26.265 106.450 26.275 ;
        RECT 106.080 26.005 107.155 26.265 ;
        RECT 108.680 26.050 110.310 26.330 ;
        RECT 111.405 26.265 111.775 26.275 ;
        RECT 111.405 26.005 112.480 26.265 ;
        RECT 114.005 26.050 115.635 26.330 ;
        RECT 116.740 26.265 117.110 26.275 ;
        RECT 116.740 26.005 117.815 26.265 ;
        RECT 119.340 26.050 120.970 26.330 ;
        RECT 36.785 25.995 37.155 26.005 ;
        RECT 42.120 25.995 42.490 26.005 ;
        RECT 47.445 25.995 47.815 26.005 ;
        RECT 52.780 25.995 53.150 26.005 ;
        RECT 58.105 25.995 58.475 26.005 ;
        RECT 63.440 25.995 63.810 26.005 ;
        RECT 68.765 25.995 69.135 26.005 ;
        RECT 74.100 25.995 74.470 26.005 ;
        RECT 79.425 25.995 79.795 26.005 ;
        RECT 84.760 25.995 85.130 26.005 ;
        RECT 90.085 25.995 90.455 26.005 ;
        RECT 95.420 25.995 95.790 26.005 ;
        RECT 100.745 25.995 101.115 26.005 ;
        RECT 106.080 25.995 106.450 26.005 ;
        RECT 111.405 25.995 111.775 26.005 ;
        RECT 116.740 25.995 117.110 26.005 ;
        RECT 41.290 25.635 41.660 25.645 ;
        RECT 46.625 25.635 46.995 25.645 ;
        RECT 51.950 25.635 52.320 25.645 ;
        RECT 57.285 25.635 57.655 25.645 ;
        RECT 62.610 25.635 62.980 25.645 ;
        RECT 67.945 25.635 68.315 25.645 ;
        RECT 73.270 25.635 73.640 25.645 ;
        RECT 78.605 25.635 78.975 25.645 ;
        RECT 83.930 25.635 84.300 25.645 ;
        RECT 89.265 25.635 89.635 25.645 ;
        RECT 94.590 25.635 94.960 25.645 ;
        RECT 99.925 25.635 100.295 25.645 ;
        RECT 105.250 25.635 105.620 25.645 ;
        RECT 110.585 25.635 110.955 25.645 ;
        RECT 115.910 25.635 116.280 25.645 ;
        RECT 121.245 25.635 121.615 25.645 ;
        RECT 40.630 25.375 41.660 25.635 ;
        RECT 45.965 25.375 46.995 25.635 ;
        RECT 51.290 25.375 52.320 25.635 ;
        RECT 56.625 25.375 57.655 25.635 ;
        RECT 61.950 25.375 62.980 25.635 ;
        RECT 67.285 25.375 68.315 25.635 ;
        RECT 72.610 25.375 73.640 25.635 ;
        RECT 77.945 25.375 78.975 25.635 ;
        RECT 83.270 25.375 84.300 25.635 ;
        RECT 88.605 25.375 89.635 25.635 ;
        RECT 93.930 25.375 94.960 25.635 ;
        RECT 99.265 25.375 100.295 25.635 ;
        RECT 104.590 25.375 105.620 25.635 ;
        RECT 109.925 25.375 110.955 25.635 ;
        RECT 115.250 25.375 116.280 25.635 ;
        RECT 120.585 25.375 121.615 25.635 ;
        RECT 41.290 25.365 41.660 25.375 ;
        RECT 46.625 25.365 46.995 25.375 ;
        RECT 51.950 25.365 52.320 25.375 ;
        RECT 57.285 25.365 57.655 25.375 ;
        RECT 62.610 25.365 62.980 25.375 ;
        RECT 67.945 25.365 68.315 25.375 ;
        RECT 73.270 25.365 73.640 25.375 ;
        RECT 78.605 25.365 78.975 25.375 ;
        RECT 83.930 25.365 84.300 25.375 ;
        RECT 89.265 25.365 89.635 25.375 ;
        RECT 94.590 25.365 94.960 25.375 ;
        RECT 99.925 25.365 100.295 25.375 ;
        RECT 105.250 25.365 105.620 25.375 ;
        RECT 110.585 25.365 110.955 25.375 ;
        RECT 115.910 25.365 116.280 25.375 ;
        RECT 121.245 25.365 121.615 25.375 ;
        RECT 36.790 23.900 37.160 23.910 ;
        RECT 42.125 23.900 42.495 23.910 ;
        RECT 47.450 23.900 47.820 23.910 ;
        RECT 52.785 23.900 53.155 23.910 ;
        RECT 58.110 23.900 58.480 23.910 ;
        RECT 63.445 23.900 63.815 23.910 ;
        RECT 68.770 23.900 69.140 23.910 ;
        RECT 74.105 23.900 74.475 23.910 ;
        RECT 79.430 23.900 79.800 23.910 ;
        RECT 84.765 23.900 85.135 23.910 ;
        RECT 90.090 23.900 90.460 23.910 ;
        RECT 95.425 23.900 95.795 23.910 ;
        RECT 100.750 23.900 101.120 23.910 ;
        RECT 106.085 23.900 106.455 23.910 ;
        RECT 111.410 23.900 111.780 23.910 ;
        RECT 116.745 23.900 117.115 23.910 ;
        RECT 36.790 23.640 37.810 23.900 ;
        RECT 42.125 23.640 43.145 23.900 ;
        RECT 47.450 23.640 48.470 23.900 ;
        RECT 52.785 23.640 53.805 23.900 ;
        RECT 58.110 23.640 59.130 23.900 ;
        RECT 63.445 23.640 64.465 23.900 ;
        RECT 68.770 23.640 69.790 23.900 ;
        RECT 74.105 23.640 75.125 23.900 ;
        RECT 79.430 23.640 80.450 23.900 ;
        RECT 84.765 23.640 85.785 23.900 ;
        RECT 90.090 23.640 91.110 23.900 ;
        RECT 95.425 23.640 96.445 23.900 ;
        RECT 100.750 23.640 101.770 23.900 ;
        RECT 106.085 23.640 107.105 23.900 ;
        RECT 111.410 23.640 112.430 23.900 ;
        RECT 116.745 23.640 117.765 23.900 ;
        RECT 36.790 23.630 37.160 23.640 ;
        RECT 42.125 23.630 42.495 23.640 ;
        RECT 47.450 23.630 47.820 23.640 ;
        RECT 52.785 23.630 53.155 23.640 ;
        RECT 58.110 23.630 58.480 23.640 ;
        RECT 63.445 23.630 63.815 23.640 ;
        RECT 68.770 23.630 69.140 23.640 ;
        RECT 74.105 23.630 74.475 23.640 ;
        RECT 79.430 23.630 79.800 23.640 ;
        RECT 84.765 23.630 85.135 23.640 ;
        RECT 90.090 23.630 90.460 23.640 ;
        RECT 95.425 23.630 95.795 23.640 ;
        RECT 100.750 23.630 101.120 23.640 ;
        RECT 106.085 23.630 106.455 23.640 ;
        RECT 111.410 23.630 111.780 23.640 ;
        RECT 116.745 23.630 117.115 23.640 ;
        RECT 41.285 23.250 41.655 23.260 ;
        RECT 46.620 23.250 46.990 23.260 ;
        RECT 51.945 23.250 52.315 23.260 ;
        RECT 57.280 23.250 57.650 23.260 ;
        RECT 62.605 23.250 62.975 23.260 ;
        RECT 67.940 23.250 68.310 23.260 ;
        RECT 73.265 23.250 73.635 23.260 ;
        RECT 78.600 23.250 78.970 23.260 ;
        RECT 83.925 23.250 84.295 23.260 ;
        RECT 89.260 23.250 89.630 23.260 ;
        RECT 94.585 23.250 94.955 23.260 ;
        RECT 99.920 23.250 100.290 23.260 ;
        RECT 105.245 23.250 105.615 23.260 ;
        RECT 110.580 23.250 110.950 23.260 ;
        RECT 115.905 23.250 116.275 23.260 ;
        RECT 121.240 23.250 121.610 23.260 ;
        RECT 37.430 22.775 39.055 23.055 ;
        RECT 40.580 22.990 41.655 23.250 ;
        RECT 41.285 22.980 41.655 22.990 ;
        RECT 42.765 22.775 44.390 23.055 ;
        RECT 45.915 22.990 46.990 23.250 ;
        RECT 46.620 22.980 46.990 22.990 ;
        RECT 48.090 22.775 49.715 23.055 ;
        RECT 51.240 22.990 52.315 23.250 ;
        RECT 51.945 22.980 52.315 22.990 ;
        RECT 53.425 22.775 55.050 23.055 ;
        RECT 56.575 22.990 57.650 23.250 ;
        RECT 57.280 22.980 57.650 22.990 ;
        RECT 58.750 22.775 60.375 23.055 ;
        RECT 61.900 22.990 62.975 23.250 ;
        RECT 62.605 22.980 62.975 22.990 ;
        RECT 64.085 22.775 65.710 23.055 ;
        RECT 67.235 22.990 68.310 23.250 ;
        RECT 67.940 22.980 68.310 22.990 ;
        RECT 69.410 22.775 71.035 23.055 ;
        RECT 72.560 22.990 73.635 23.250 ;
        RECT 73.265 22.980 73.635 22.990 ;
        RECT 74.745 22.775 76.370 23.055 ;
        RECT 77.895 22.990 78.970 23.250 ;
        RECT 78.600 22.980 78.970 22.990 ;
        RECT 80.070 22.775 81.695 23.055 ;
        RECT 83.220 22.990 84.295 23.250 ;
        RECT 83.925 22.980 84.295 22.990 ;
        RECT 85.405 22.775 87.030 23.055 ;
        RECT 88.555 22.990 89.630 23.250 ;
        RECT 89.260 22.980 89.630 22.990 ;
        RECT 90.730 22.775 92.355 23.055 ;
        RECT 93.880 22.990 94.955 23.250 ;
        RECT 94.585 22.980 94.955 22.990 ;
        RECT 96.065 22.775 97.690 23.055 ;
        RECT 99.215 22.990 100.290 23.250 ;
        RECT 99.920 22.980 100.290 22.990 ;
        RECT 101.390 22.775 103.015 23.055 ;
        RECT 104.540 22.990 105.615 23.250 ;
        RECT 105.245 22.980 105.615 22.990 ;
        RECT 106.725 22.775 108.350 23.055 ;
        RECT 109.875 22.990 110.950 23.250 ;
        RECT 110.580 22.980 110.950 22.990 ;
        RECT 112.050 22.775 113.675 23.055 ;
        RECT 115.200 22.990 116.275 23.250 ;
        RECT 115.905 22.980 116.275 22.990 ;
        RECT 117.385 22.775 119.010 23.055 ;
        RECT 120.535 22.990 121.610 23.250 ;
        RECT 121.240 22.980 121.610 22.990 ;
        RECT 38.795 22.555 39.055 22.775 ;
        RECT 44.130 22.555 44.390 22.775 ;
        RECT 49.455 22.555 49.715 22.775 ;
        RECT 54.790 22.555 55.050 22.775 ;
        RECT 60.115 22.555 60.375 22.775 ;
        RECT 65.450 22.555 65.710 22.775 ;
        RECT 70.775 22.555 71.035 22.775 ;
        RECT 76.110 22.555 76.370 22.775 ;
        RECT 81.435 22.555 81.695 22.775 ;
        RECT 86.770 22.555 87.030 22.775 ;
        RECT 92.095 22.555 92.355 22.775 ;
        RECT 97.430 22.555 97.690 22.775 ;
        RECT 102.755 22.555 103.015 22.775 ;
        RECT 108.090 22.555 108.350 22.775 ;
        RECT 113.415 22.555 113.675 22.775 ;
        RECT 118.750 22.555 119.010 22.775 ;
        RECT 32.625 22.275 34.390 22.555 ;
        RECT 37.950 22.275 38.470 22.555 ;
        RECT 38.715 22.275 39.110 22.555 ;
        RECT 39.330 22.275 39.730 22.555 ;
        RECT 43.285 22.275 43.805 22.555 ;
        RECT 44.050 22.275 44.445 22.555 ;
        RECT 44.665 22.275 45.065 22.555 ;
        RECT 48.610 22.275 49.130 22.555 ;
        RECT 49.375 22.275 49.770 22.555 ;
        RECT 49.990 22.275 50.390 22.555 ;
        RECT 53.945 22.275 54.465 22.555 ;
        RECT 54.710 22.275 55.105 22.555 ;
        RECT 55.325 22.275 55.725 22.555 ;
        RECT 59.270 22.275 59.790 22.555 ;
        RECT 60.035 22.275 60.430 22.555 ;
        RECT 60.650 22.275 61.050 22.555 ;
        RECT 64.605 22.275 65.125 22.555 ;
        RECT 65.370 22.275 65.765 22.555 ;
        RECT 65.985 22.275 66.385 22.555 ;
        RECT 69.930 22.275 70.450 22.555 ;
        RECT 70.695 22.275 71.090 22.555 ;
        RECT 71.310 22.275 71.710 22.555 ;
        RECT 75.265 22.275 75.785 22.555 ;
        RECT 76.030 22.275 76.425 22.555 ;
        RECT 76.645 22.275 77.045 22.555 ;
        RECT 80.590 22.275 81.110 22.555 ;
        RECT 81.355 22.275 81.750 22.555 ;
        RECT 81.970 22.275 82.370 22.555 ;
        RECT 85.925 22.275 86.445 22.555 ;
        RECT 86.690 22.275 87.085 22.555 ;
        RECT 87.305 22.275 87.705 22.555 ;
        RECT 91.250 22.275 91.770 22.555 ;
        RECT 92.015 22.275 92.410 22.555 ;
        RECT 92.630 22.275 93.030 22.555 ;
        RECT 96.585 22.275 97.105 22.555 ;
        RECT 97.350 22.275 97.745 22.555 ;
        RECT 97.965 22.275 98.365 22.555 ;
        RECT 101.910 22.275 102.430 22.555 ;
        RECT 102.675 22.275 103.070 22.555 ;
        RECT 103.290 22.275 103.690 22.555 ;
        RECT 107.245 22.275 107.765 22.555 ;
        RECT 108.010 22.275 108.405 22.555 ;
        RECT 108.625 22.275 109.025 22.555 ;
        RECT 112.570 22.275 113.090 22.555 ;
        RECT 113.335 22.275 113.730 22.555 ;
        RECT 113.950 22.275 114.350 22.555 ;
        RECT 117.905 22.275 118.425 22.555 ;
        RECT 118.670 22.275 119.065 22.555 ;
        RECT 119.285 22.275 119.685 22.555 ;
        RECT 123.230 22.275 124.995 22.555 ;
        RECT 36.785 22.055 37.155 22.065 ;
        RECT 42.120 22.055 42.490 22.065 ;
        RECT 47.445 22.055 47.815 22.065 ;
        RECT 52.780 22.055 53.150 22.065 ;
        RECT 58.105 22.055 58.475 22.065 ;
        RECT 63.440 22.055 63.810 22.065 ;
        RECT 68.765 22.055 69.135 22.065 ;
        RECT 74.100 22.055 74.470 22.065 ;
        RECT 79.425 22.055 79.795 22.065 ;
        RECT 84.760 22.055 85.130 22.065 ;
        RECT 90.085 22.055 90.455 22.065 ;
        RECT 95.420 22.055 95.790 22.065 ;
        RECT 100.745 22.055 101.115 22.065 ;
        RECT 106.080 22.055 106.450 22.065 ;
        RECT 111.405 22.055 111.775 22.065 ;
        RECT 116.740 22.055 117.110 22.065 ;
        RECT 36.785 21.795 37.810 22.055 ;
        RECT 41.285 21.965 41.655 21.975 ;
        RECT 36.785 21.785 37.155 21.795 ;
        RECT 28.415 21.345 28.695 21.715 ;
        RECT 40.630 21.705 41.655 21.965 ;
        RECT 42.120 21.795 43.145 22.055 ;
        RECT 46.620 21.965 46.990 21.975 ;
        RECT 42.120 21.785 42.490 21.795 ;
        RECT 45.965 21.705 46.990 21.965 ;
        RECT 47.445 21.795 48.470 22.055 ;
        RECT 51.945 21.965 52.315 21.975 ;
        RECT 47.445 21.785 47.815 21.795 ;
        RECT 51.290 21.705 52.315 21.965 ;
        RECT 52.780 21.795 53.805 22.055 ;
        RECT 57.280 21.965 57.650 21.975 ;
        RECT 52.780 21.785 53.150 21.795 ;
        RECT 56.625 21.705 57.650 21.965 ;
        RECT 58.105 21.795 59.130 22.055 ;
        RECT 62.605 21.965 62.975 21.975 ;
        RECT 58.105 21.785 58.475 21.795 ;
        RECT 61.950 21.705 62.975 21.965 ;
        RECT 63.440 21.795 64.465 22.055 ;
        RECT 67.940 21.965 68.310 21.975 ;
        RECT 63.440 21.785 63.810 21.795 ;
        RECT 67.285 21.705 68.310 21.965 ;
        RECT 68.765 21.795 69.790 22.055 ;
        RECT 73.265 21.965 73.635 21.975 ;
        RECT 68.765 21.785 69.135 21.795 ;
        RECT 72.610 21.705 73.635 21.965 ;
        RECT 74.100 21.795 75.125 22.055 ;
        RECT 78.600 21.965 78.970 21.975 ;
        RECT 74.100 21.785 74.470 21.795 ;
        RECT 77.945 21.705 78.970 21.965 ;
        RECT 79.425 21.795 80.450 22.055 ;
        RECT 83.925 21.965 84.295 21.975 ;
        RECT 79.425 21.785 79.795 21.795 ;
        RECT 83.270 21.705 84.295 21.965 ;
        RECT 84.760 21.795 85.785 22.055 ;
        RECT 89.260 21.965 89.630 21.975 ;
        RECT 84.760 21.785 85.130 21.795 ;
        RECT 88.605 21.705 89.630 21.965 ;
        RECT 90.085 21.795 91.110 22.055 ;
        RECT 94.585 21.965 94.955 21.975 ;
        RECT 90.085 21.785 90.455 21.795 ;
        RECT 93.930 21.705 94.955 21.965 ;
        RECT 95.420 21.795 96.445 22.055 ;
        RECT 99.920 21.965 100.290 21.975 ;
        RECT 95.420 21.785 95.790 21.795 ;
        RECT 99.265 21.705 100.290 21.965 ;
        RECT 100.745 21.795 101.770 22.055 ;
        RECT 105.245 21.965 105.615 21.975 ;
        RECT 100.745 21.785 101.115 21.795 ;
        RECT 104.590 21.705 105.615 21.965 ;
        RECT 106.080 21.795 107.105 22.055 ;
        RECT 110.580 21.965 110.950 21.975 ;
        RECT 106.080 21.785 106.450 21.795 ;
        RECT 109.925 21.705 110.950 21.965 ;
        RECT 111.405 21.795 112.430 22.055 ;
        RECT 115.905 21.965 116.275 21.975 ;
        RECT 111.405 21.785 111.775 21.795 ;
        RECT 115.250 21.705 116.275 21.965 ;
        RECT 116.740 21.795 117.765 22.055 ;
        RECT 121.240 21.965 121.610 21.975 ;
        RECT 116.740 21.785 117.110 21.795 ;
        RECT 120.585 21.705 121.610 21.965 ;
        RECT 41.285 21.695 41.655 21.705 ;
        RECT 46.620 21.695 46.990 21.705 ;
        RECT 51.945 21.695 52.315 21.705 ;
        RECT 57.280 21.695 57.650 21.705 ;
        RECT 62.605 21.695 62.975 21.705 ;
        RECT 67.940 21.695 68.310 21.705 ;
        RECT 73.265 21.695 73.635 21.705 ;
        RECT 78.600 21.695 78.970 21.705 ;
        RECT 83.925 21.695 84.295 21.705 ;
        RECT 89.260 21.695 89.630 21.705 ;
        RECT 94.585 21.695 94.955 21.705 ;
        RECT 99.920 21.695 100.290 21.705 ;
        RECT 105.245 21.695 105.615 21.705 ;
        RECT 110.580 21.695 110.950 21.705 ;
        RECT 115.905 21.695 116.275 21.705 ;
        RECT 121.240 21.695 121.610 21.705 ;
        RECT 28.030 20.015 28.310 20.385 ;
        RECT 27.655 19.365 27.935 19.735 ;
        RECT 27.275 18.075 27.555 18.445 ;
        RECT 27.325 14.825 27.505 18.075 ;
        RECT 27.705 17.475 27.885 19.365 ;
        RECT 27.665 16.370 27.925 17.475 ;
        RECT 27.705 16.115 27.885 16.370 ;
        RECT 27.650 15.745 27.930 16.115 ;
        RECT 27.705 15.695 27.885 15.745 ;
        RECT 27.275 14.455 27.555 14.825 ;
        RECT 27.325 12.150 27.505 14.455 ;
        RECT 28.085 14.180 28.265 20.015 ;
        RECT 28.465 19.090 28.645 21.345 ;
        RECT 36.785 20.030 37.155 20.040 ;
        RECT 42.120 20.030 42.490 20.040 ;
        RECT 47.445 20.030 47.815 20.040 ;
        RECT 52.780 20.030 53.150 20.040 ;
        RECT 58.105 20.030 58.475 20.040 ;
        RECT 63.440 20.030 63.810 20.040 ;
        RECT 68.765 20.030 69.135 20.040 ;
        RECT 74.100 20.030 74.470 20.040 ;
        RECT 79.425 20.030 79.795 20.040 ;
        RECT 84.760 20.030 85.130 20.040 ;
        RECT 90.085 20.030 90.455 20.040 ;
        RECT 95.420 20.030 95.790 20.040 ;
        RECT 100.745 20.030 101.115 20.040 ;
        RECT 106.080 20.030 106.450 20.040 ;
        RECT 111.405 20.030 111.775 20.040 ;
        RECT 116.740 20.030 117.110 20.040 ;
        RECT 36.785 19.770 37.810 20.030 ;
        RECT 41.285 19.935 41.655 19.945 ;
        RECT 36.785 19.760 37.155 19.770 ;
        RECT 40.630 19.675 41.655 19.935 ;
        RECT 42.120 19.770 43.145 20.030 ;
        RECT 46.620 19.935 46.990 19.945 ;
        RECT 42.120 19.760 42.490 19.770 ;
        RECT 45.965 19.675 46.990 19.935 ;
        RECT 47.445 19.770 48.470 20.030 ;
        RECT 51.945 19.935 52.315 19.945 ;
        RECT 47.445 19.760 47.815 19.770 ;
        RECT 51.290 19.675 52.315 19.935 ;
        RECT 52.780 19.770 53.805 20.030 ;
        RECT 57.280 19.935 57.650 19.945 ;
        RECT 52.780 19.760 53.150 19.770 ;
        RECT 56.625 19.675 57.650 19.935 ;
        RECT 58.105 19.770 59.130 20.030 ;
        RECT 62.605 19.935 62.975 19.945 ;
        RECT 58.105 19.760 58.475 19.770 ;
        RECT 61.950 19.675 62.975 19.935 ;
        RECT 63.440 19.770 64.465 20.030 ;
        RECT 67.940 19.935 68.310 19.945 ;
        RECT 63.440 19.760 63.810 19.770 ;
        RECT 67.285 19.675 68.310 19.935 ;
        RECT 68.765 19.770 69.790 20.030 ;
        RECT 73.265 19.935 73.635 19.945 ;
        RECT 68.765 19.760 69.135 19.770 ;
        RECT 72.610 19.675 73.635 19.935 ;
        RECT 74.100 19.770 75.125 20.030 ;
        RECT 78.600 19.935 78.970 19.945 ;
        RECT 74.100 19.760 74.470 19.770 ;
        RECT 77.945 19.675 78.970 19.935 ;
        RECT 79.425 19.770 80.450 20.030 ;
        RECT 83.925 19.935 84.295 19.945 ;
        RECT 79.425 19.760 79.795 19.770 ;
        RECT 83.270 19.675 84.295 19.935 ;
        RECT 84.760 19.770 85.785 20.030 ;
        RECT 89.260 19.935 89.630 19.945 ;
        RECT 84.760 19.760 85.130 19.770 ;
        RECT 88.605 19.675 89.630 19.935 ;
        RECT 90.085 19.770 91.110 20.030 ;
        RECT 94.585 19.935 94.955 19.945 ;
        RECT 90.085 19.760 90.455 19.770 ;
        RECT 93.930 19.675 94.955 19.935 ;
        RECT 95.420 19.770 96.445 20.030 ;
        RECT 99.920 19.935 100.290 19.945 ;
        RECT 95.420 19.760 95.790 19.770 ;
        RECT 99.265 19.675 100.290 19.935 ;
        RECT 100.745 19.770 101.770 20.030 ;
        RECT 105.245 19.935 105.615 19.945 ;
        RECT 100.745 19.760 101.115 19.770 ;
        RECT 104.590 19.675 105.615 19.935 ;
        RECT 106.080 19.770 107.105 20.030 ;
        RECT 110.580 19.935 110.950 19.945 ;
        RECT 106.080 19.760 106.450 19.770 ;
        RECT 109.925 19.675 110.950 19.935 ;
        RECT 111.405 19.770 112.430 20.030 ;
        RECT 115.905 19.935 116.275 19.945 ;
        RECT 111.405 19.760 111.775 19.770 ;
        RECT 115.250 19.675 116.275 19.935 ;
        RECT 116.740 19.770 117.765 20.030 ;
        RECT 121.240 19.935 121.610 19.945 ;
        RECT 116.740 19.760 117.110 19.770 ;
        RECT 120.585 19.675 121.610 19.935 ;
        RECT 41.285 19.665 41.655 19.675 ;
        RECT 46.620 19.665 46.990 19.675 ;
        RECT 51.945 19.665 52.315 19.675 ;
        RECT 57.280 19.665 57.650 19.675 ;
        RECT 62.605 19.665 62.975 19.675 ;
        RECT 67.940 19.665 68.310 19.675 ;
        RECT 73.265 19.665 73.635 19.675 ;
        RECT 78.600 19.665 78.970 19.675 ;
        RECT 83.925 19.665 84.295 19.675 ;
        RECT 89.260 19.665 89.630 19.675 ;
        RECT 94.585 19.665 94.955 19.675 ;
        RECT 99.920 19.665 100.290 19.675 ;
        RECT 105.245 19.665 105.615 19.675 ;
        RECT 110.580 19.665 110.950 19.675 ;
        RECT 115.905 19.665 116.275 19.675 ;
        RECT 121.240 19.665 121.610 19.675 ;
        RECT 34.005 19.380 34.400 19.385 ;
        RECT 33.390 19.100 35.160 19.380 ;
        RECT 38.715 19.100 39.110 19.380 ;
        RECT 39.330 19.105 39.730 19.385 ;
        RECT 40.120 19.100 41.025 19.380 ;
        RECT 44.050 19.100 44.445 19.380 ;
        RECT 44.665 19.105 45.065 19.385 ;
        RECT 45.455 19.100 46.360 19.380 ;
        RECT 49.375 19.100 49.770 19.380 ;
        RECT 49.990 19.105 50.390 19.385 ;
        RECT 50.780 19.100 51.685 19.380 ;
        RECT 54.710 19.100 55.105 19.380 ;
        RECT 55.325 19.105 55.725 19.385 ;
        RECT 56.115 19.100 57.020 19.380 ;
        RECT 60.035 19.100 60.430 19.380 ;
        RECT 60.650 19.105 61.050 19.385 ;
        RECT 61.440 19.100 62.345 19.380 ;
        RECT 65.370 19.100 65.765 19.380 ;
        RECT 65.985 19.105 66.385 19.385 ;
        RECT 66.775 19.100 67.680 19.380 ;
        RECT 70.695 19.100 71.090 19.380 ;
        RECT 71.310 19.105 71.710 19.385 ;
        RECT 72.100 19.100 73.005 19.380 ;
        RECT 76.030 19.100 76.425 19.380 ;
        RECT 76.645 19.105 77.045 19.385 ;
        RECT 77.435 19.100 78.340 19.380 ;
        RECT 81.355 19.100 81.750 19.380 ;
        RECT 81.970 19.105 82.370 19.385 ;
        RECT 82.760 19.100 83.665 19.380 ;
        RECT 86.690 19.100 87.085 19.380 ;
        RECT 87.305 19.105 87.705 19.385 ;
        RECT 88.095 19.100 89.000 19.380 ;
        RECT 92.015 19.100 92.410 19.380 ;
        RECT 92.630 19.105 93.030 19.385 ;
        RECT 93.420 19.100 94.325 19.380 ;
        RECT 97.350 19.100 97.745 19.380 ;
        RECT 97.965 19.105 98.365 19.385 ;
        RECT 98.755 19.100 99.660 19.380 ;
        RECT 102.675 19.100 103.070 19.380 ;
        RECT 103.290 19.105 103.690 19.385 ;
        RECT 104.080 19.100 104.985 19.380 ;
        RECT 108.010 19.100 108.405 19.380 ;
        RECT 108.625 19.105 109.025 19.385 ;
        RECT 109.415 19.100 110.320 19.380 ;
        RECT 113.335 19.100 113.730 19.380 ;
        RECT 113.950 19.105 114.350 19.385 ;
        RECT 114.740 19.100 115.645 19.380 ;
        RECT 118.670 19.100 119.065 19.380 ;
        RECT 119.285 19.105 119.685 19.385 ;
        RECT 124.610 19.380 125.005 19.385 ;
        RECT 120.075 19.100 120.980 19.380 ;
        RECT 123.995 19.100 125.765 19.380 ;
        RECT 28.415 18.720 28.695 19.090 ;
        RECT 36.785 18.730 37.155 18.740 ;
        RECT 42.120 18.730 42.490 18.740 ;
        RECT 47.445 18.730 47.815 18.740 ;
        RECT 52.780 18.730 53.150 18.740 ;
        RECT 58.105 18.730 58.475 18.740 ;
        RECT 63.440 18.730 63.810 18.740 ;
        RECT 68.765 18.730 69.135 18.740 ;
        RECT 74.100 18.730 74.470 18.740 ;
        RECT 79.425 18.730 79.795 18.740 ;
        RECT 84.760 18.730 85.130 18.740 ;
        RECT 90.085 18.730 90.455 18.740 ;
        RECT 95.420 18.730 95.790 18.740 ;
        RECT 100.745 18.730 101.115 18.740 ;
        RECT 106.080 18.730 106.450 18.740 ;
        RECT 111.405 18.730 111.775 18.740 ;
        RECT 116.740 18.730 117.110 18.740 ;
        RECT 28.465 15.470 28.645 18.720 ;
        RECT 36.785 18.470 37.860 18.730 ;
        RECT 42.120 18.470 43.195 18.730 ;
        RECT 47.445 18.470 48.520 18.730 ;
        RECT 52.780 18.470 53.855 18.730 ;
        RECT 58.105 18.470 59.180 18.730 ;
        RECT 63.440 18.470 64.515 18.730 ;
        RECT 68.765 18.470 69.840 18.730 ;
        RECT 74.100 18.470 75.175 18.730 ;
        RECT 79.425 18.470 80.500 18.730 ;
        RECT 84.760 18.470 85.835 18.730 ;
        RECT 90.085 18.470 91.160 18.730 ;
        RECT 95.420 18.470 96.495 18.730 ;
        RECT 100.745 18.470 101.820 18.730 ;
        RECT 106.080 18.470 107.155 18.730 ;
        RECT 111.405 18.470 112.480 18.730 ;
        RECT 116.740 18.470 117.815 18.730 ;
        RECT 36.785 18.460 37.155 18.470 ;
        RECT 42.120 18.460 42.490 18.470 ;
        RECT 47.445 18.460 47.815 18.470 ;
        RECT 52.780 18.460 53.150 18.470 ;
        RECT 58.105 18.460 58.475 18.470 ;
        RECT 63.440 18.460 63.810 18.470 ;
        RECT 68.765 18.460 69.135 18.470 ;
        RECT 74.100 18.460 74.470 18.470 ;
        RECT 79.425 18.460 79.795 18.470 ;
        RECT 84.760 18.460 85.130 18.470 ;
        RECT 90.085 18.460 90.455 18.470 ;
        RECT 95.420 18.460 95.790 18.470 ;
        RECT 100.745 18.460 101.115 18.470 ;
        RECT 106.080 18.460 106.450 18.470 ;
        RECT 111.405 18.460 111.775 18.470 ;
        RECT 116.740 18.460 117.110 18.470 ;
        RECT 41.290 18.100 41.660 18.110 ;
        RECT 46.625 18.100 46.995 18.110 ;
        RECT 51.950 18.100 52.320 18.110 ;
        RECT 57.285 18.100 57.655 18.110 ;
        RECT 62.610 18.100 62.980 18.110 ;
        RECT 67.945 18.100 68.315 18.110 ;
        RECT 73.270 18.100 73.640 18.110 ;
        RECT 78.605 18.100 78.975 18.110 ;
        RECT 83.930 18.100 84.300 18.110 ;
        RECT 89.265 18.100 89.635 18.110 ;
        RECT 94.590 18.100 94.960 18.110 ;
        RECT 99.925 18.100 100.295 18.110 ;
        RECT 105.250 18.100 105.620 18.110 ;
        RECT 110.585 18.100 110.955 18.110 ;
        RECT 115.910 18.100 116.280 18.110 ;
        RECT 121.245 18.100 121.615 18.110 ;
        RECT 40.630 17.840 41.660 18.100 ;
        RECT 45.965 17.840 46.995 18.100 ;
        RECT 51.290 17.840 52.320 18.100 ;
        RECT 56.625 17.840 57.655 18.100 ;
        RECT 61.950 17.840 62.980 18.100 ;
        RECT 67.285 17.840 68.315 18.100 ;
        RECT 72.610 17.840 73.640 18.100 ;
        RECT 77.945 17.840 78.975 18.100 ;
        RECT 83.270 17.840 84.300 18.100 ;
        RECT 88.605 17.840 89.635 18.100 ;
        RECT 93.930 17.840 94.960 18.100 ;
        RECT 99.265 17.840 100.295 18.100 ;
        RECT 104.590 17.840 105.620 18.100 ;
        RECT 109.925 17.840 110.955 18.100 ;
        RECT 115.250 17.840 116.280 18.100 ;
        RECT 120.585 17.840 121.615 18.100 ;
        RECT 41.290 17.830 41.660 17.840 ;
        RECT 46.625 17.830 46.995 17.840 ;
        RECT 51.950 17.830 52.320 17.840 ;
        RECT 57.285 17.830 57.655 17.840 ;
        RECT 62.610 17.830 62.980 17.840 ;
        RECT 67.945 17.830 68.315 17.840 ;
        RECT 73.270 17.830 73.640 17.840 ;
        RECT 78.605 17.830 78.975 17.840 ;
        RECT 83.930 17.830 84.300 17.840 ;
        RECT 89.265 17.830 89.635 17.840 ;
        RECT 94.590 17.830 94.960 17.840 ;
        RECT 99.925 17.830 100.295 17.840 ;
        RECT 105.250 17.830 105.620 17.840 ;
        RECT 110.585 17.830 110.955 17.840 ;
        RECT 115.910 17.830 116.280 17.840 ;
        RECT 121.245 17.830 121.615 17.840 ;
        RECT 36.790 16.365 37.160 16.375 ;
        RECT 42.125 16.365 42.495 16.375 ;
        RECT 47.450 16.365 47.820 16.375 ;
        RECT 52.785 16.365 53.155 16.375 ;
        RECT 58.110 16.365 58.480 16.375 ;
        RECT 63.445 16.365 63.815 16.375 ;
        RECT 68.770 16.365 69.140 16.375 ;
        RECT 74.105 16.365 74.475 16.375 ;
        RECT 79.430 16.365 79.800 16.375 ;
        RECT 84.765 16.365 85.135 16.375 ;
        RECT 90.090 16.365 90.460 16.375 ;
        RECT 95.425 16.365 95.795 16.375 ;
        RECT 100.750 16.365 101.120 16.375 ;
        RECT 106.085 16.365 106.455 16.375 ;
        RECT 111.410 16.365 111.780 16.375 ;
        RECT 116.745 16.365 117.115 16.375 ;
        RECT 36.790 16.105 37.810 16.365 ;
        RECT 42.125 16.105 43.145 16.365 ;
        RECT 47.450 16.105 48.470 16.365 ;
        RECT 52.785 16.105 53.805 16.365 ;
        RECT 58.110 16.105 59.130 16.365 ;
        RECT 63.445 16.105 64.465 16.365 ;
        RECT 68.770 16.105 69.790 16.365 ;
        RECT 74.105 16.105 75.125 16.365 ;
        RECT 79.430 16.105 80.450 16.365 ;
        RECT 84.765 16.105 85.785 16.365 ;
        RECT 90.090 16.105 91.110 16.365 ;
        RECT 95.425 16.105 96.445 16.365 ;
        RECT 100.750 16.105 101.770 16.365 ;
        RECT 106.085 16.105 107.105 16.365 ;
        RECT 111.410 16.105 112.430 16.365 ;
        RECT 116.745 16.105 117.765 16.365 ;
        RECT 36.790 16.095 37.160 16.105 ;
        RECT 42.125 16.095 42.495 16.105 ;
        RECT 47.450 16.095 47.820 16.105 ;
        RECT 52.785 16.095 53.155 16.105 ;
        RECT 58.110 16.095 58.480 16.105 ;
        RECT 63.445 16.095 63.815 16.105 ;
        RECT 68.770 16.095 69.140 16.105 ;
        RECT 74.105 16.095 74.475 16.105 ;
        RECT 79.430 16.095 79.800 16.105 ;
        RECT 84.765 16.095 85.135 16.105 ;
        RECT 90.090 16.095 90.460 16.105 ;
        RECT 95.425 16.095 95.795 16.105 ;
        RECT 100.750 16.095 101.120 16.105 ;
        RECT 106.085 16.095 106.455 16.105 ;
        RECT 111.410 16.095 111.780 16.105 ;
        RECT 116.745 16.095 117.115 16.105 ;
        RECT 41.285 15.715 41.655 15.725 ;
        RECT 46.620 15.715 46.990 15.725 ;
        RECT 51.945 15.715 52.315 15.725 ;
        RECT 57.280 15.715 57.650 15.725 ;
        RECT 62.605 15.715 62.975 15.725 ;
        RECT 67.940 15.715 68.310 15.725 ;
        RECT 73.265 15.715 73.635 15.725 ;
        RECT 78.600 15.715 78.970 15.725 ;
        RECT 83.925 15.715 84.295 15.725 ;
        RECT 89.260 15.715 89.630 15.725 ;
        RECT 94.585 15.715 94.955 15.725 ;
        RECT 99.920 15.715 100.290 15.725 ;
        RECT 105.245 15.715 105.615 15.725 ;
        RECT 110.580 15.715 110.950 15.725 ;
        RECT 115.905 15.715 116.275 15.725 ;
        RECT 121.240 15.715 121.610 15.725 ;
        RECT 28.415 15.100 28.695 15.470 ;
        RECT 40.580 15.455 41.655 15.715 ;
        RECT 45.915 15.455 46.990 15.715 ;
        RECT 51.240 15.455 52.315 15.715 ;
        RECT 56.575 15.455 57.650 15.715 ;
        RECT 61.900 15.455 62.975 15.715 ;
        RECT 67.235 15.455 68.310 15.715 ;
        RECT 72.560 15.455 73.635 15.715 ;
        RECT 77.895 15.455 78.970 15.715 ;
        RECT 83.220 15.455 84.295 15.715 ;
        RECT 88.555 15.455 89.630 15.715 ;
        RECT 93.880 15.455 94.955 15.715 ;
        RECT 99.215 15.455 100.290 15.715 ;
        RECT 104.540 15.455 105.615 15.715 ;
        RECT 109.875 15.455 110.950 15.715 ;
        RECT 115.200 15.455 116.275 15.715 ;
        RECT 120.535 15.455 121.610 15.715 ;
        RECT 41.285 15.445 41.655 15.455 ;
        RECT 46.620 15.445 46.990 15.455 ;
        RECT 51.945 15.445 52.315 15.455 ;
        RECT 57.280 15.445 57.650 15.455 ;
        RECT 62.605 15.445 62.975 15.455 ;
        RECT 67.940 15.445 68.310 15.455 ;
        RECT 73.265 15.445 73.635 15.455 ;
        RECT 78.600 15.445 78.970 15.455 ;
        RECT 83.925 15.445 84.295 15.455 ;
        RECT 89.260 15.445 89.630 15.455 ;
        RECT 94.585 15.445 94.955 15.455 ;
        RECT 99.920 15.445 100.290 15.455 ;
        RECT 105.245 15.445 105.615 15.455 ;
        RECT 110.580 15.445 110.950 15.455 ;
        RECT 115.905 15.445 116.275 15.455 ;
        RECT 121.240 15.445 121.610 15.455 ;
        RECT 28.035 13.810 28.315 14.180 ;
        RECT 27.285 11.045 27.545 12.150 ;
        RECT 28.085 11.550 28.265 13.810 ;
        RECT 28.465 12.845 28.645 15.100 ;
        RECT 32.625 14.740 34.390 15.020 ;
        RECT 37.950 14.740 38.470 15.020 ;
        RECT 38.715 14.740 39.110 15.020 ;
        RECT 39.330 14.740 39.730 15.020 ;
        RECT 43.285 14.740 43.805 15.020 ;
        RECT 44.050 14.740 44.445 15.020 ;
        RECT 44.665 14.740 45.065 15.020 ;
        RECT 48.610 14.740 49.130 15.020 ;
        RECT 49.375 14.740 49.770 15.020 ;
        RECT 49.990 14.740 50.390 15.020 ;
        RECT 53.945 14.740 54.465 15.020 ;
        RECT 54.710 14.740 55.105 15.020 ;
        RECT 55.325 14.740 55.725 15.020 ;
        RECT 59.270 14.740 59.790 15.020 ;
        RECT 60.035 14.740 60.430 15.020 ;
        RECT 60.650 14.740 61.050 15.020 ;
        RECT 64.605 14.740 65.125 15.020 ;
        RECT 65.370 14.740 65.765 15.020 ;
        RECT 65.985 14.740 66.385 15.020 ;
        RECT 69.930 14.740 70.450 15.020 ;
        RECT 70.695 14.740 71.090 15.020 ;
        RECT 71.310 14.740 71.710 15.020 ;
        RECT 75.265 14.740 75.785 15.020 ;
        RECT 76.030 14.740 76.425 15.020 ;
        RECT 76.645 14.740 77.045 15.020 ;
        RECT 80.590 14.740 81.110 15.020 ;
        RECT 81.355 14.740 81.750 15.020 ;
        RECT 81.970 14.740 82.370 15.020 ;
        RECT 85.925 14.740 86.445 15.020 ;
        RECT 86.690 14.740 87.085 15.020 ;
        RECT 87.305 14.740 87.705 15.020 ;
        RECT 91.250 14.740 91.770 15.020 ;
        RECT 92.015 14.740 92.410 15.020 ;
        RECT 92.630 14.740 93.030 15.020 ;
        RECT 96.585 14.740 97.105 15.020 ;
        RECT 97.350 14.740 97.745 15.020 ;
        RECT 97.965 14.740 98.365 15.020 ;
        RECT 101.910 14.740 102.430 15.020 ;
        RECT 102.675 14.740 103.070 15.020 ;
        RECT 103.290 14.740 103.690 15.020 ;
        RECT 107.245 14.740 107.765 15.020 ;
        RECT 108.010 14.740 108.405 15.020 ;
        RECT 108.625 14.740 109.025 15.020 ;
        RECT 112.570 14.740 113.090 15.020 ;
        RECT 113.335 14.740 113.730 15.020 ;
        RECT 113.950 14.740 114.350 15.020 ;
        RECT 117.905 14.740 118.425 15.020 ;
        RECT 118.670 14.740 119.065 15.020 ;
        RECT 119.285 14.740 119.685 15.020 ;
        RECT 123.230 14.740 124.995 15.020 ;
        RECT 36.785 14.520 37.155 14.530 ;
        RECT 42.120 14.520 42.490 14.530 ;
        RECT 47.445 14.520 47.815 14.530 ;
        RECT 52.780 14.520 53.150 14.530 ;
        RECT 58.105 14.520 58.475 14.530 ;
        RECT 63.440 14.520 63.810 14.530 ;
        RECT 68.765 14.520 69.135 14.530 ;
        RECT 74.100 14.520 74.470 14.530 ;
        RECT 79.425 14.520 79.795 14.530 ;
        RECT 84.760 14.520 85.130 14.530 ;
        RECT 90.085 14.520 90.455 14.530 ;
        RECT 95.420 14.520 95.790 14.530 ;
        RECT 100.745 14.520 101.115 14.530 ;
        RECT 106.080 14.520 106.450 14.530 ;
        RECT 111.405 14.520 111.775 14.530 ;
        RECT 116.740 14.520 117.110 14.530 ;
        RECT 36.785 14.260 37.810 14.520 ;
        RECT 41.285 14.430 41.655 14.440 ;
        RECT 36.785 14.250 37.155 14.260 ;
        RECT 40.630 14.170 41.655 14.430 ;
        RECT 42.120 14.260 43.145 14.520 ;
        RECT 46.620 14.430 46.990 14.440 ;
        RECT 42.120 14.250 42.490 14.260 ;
        RECT 45.965 14.170 46.990 14.430 ;
        RECT 47.445 14.260 48.470 14.520 ;
        RECT 51.945 14.430 52.315 14.440 ;
        RECT 47.445 14.250 47.815 14.260 ;
        RECT 51.290 14.170 52.315 14.430 ;
        RECT 52.780 14.260 53.805 14.520 ;
        RECT 57.280 14.430 57.650 14.440 ;
        RECT 52.780 14.250 53.150 14.260 ;
        RECT 56.625 14.170 57.650 14.430 ;
        RECT 58.105 14.260 59.130 14.520 ;
        RECT 62.605 14.430 62.975 14.440 ;
        RECT 58.105 14.250 58.475 14.260 ;
        RECT 61.950 14.170 62.975 14.430 ;
        RECT 63.440 14.260 64.465 14.520 ;
        RECT 67.940 14.430 68.310 14.440 ;
        RECT 63.440 14.250 63.810 14.260 ;
        RECT 67.285 14.170 68.310 14.430 ;
        RECT 68.765 14.260 69.790 14.520 ;
        RECT 73.265 14.430 73.635 14.440 ;
        RECT 68.765 14.250 69.135 14.260 ;
        RECT 72.610 14.170 73.635 14.430 ;
        RECT 74.100 14.260 75.125 14.520 ;
        RECT 78.600 14.430 78.970 14.440 ;
        RECT 74.100 14.250 74.470 14.260 ;
        RECT 77.945 14.170 78.970 14.430 ;
        RECT 79.425 14.260 80.450 14.520 ;
        RECT 83.925 14.430 84.295 14.440 ;
        RECT 79.425 14.250 79.795 14.260 ;
        RECT 83.270 14.170 84.295 14.430 ;
        RECT 84.760 14.260 85.785 14.520 ;
        RECT 89.260 14.430 89.630 14.440 ;
        RECT 84.760 14.250 85.130 14.260 ;
        RECT 88.605 14.170 89.630 14.430 ;
        RECT 90.085 14.260 91.110 14.520 ;
        RECT 94.585 14.430 94.955 14.440 ;
        RECT 90.085 14.250 90.455 14.260 ;
        RECT 93.930 14.170 94.955 14.430 ;
        RECT 95.420 14.260 96.445 14.520 ;
        RECT 99.920 14.430 100.290 14.440 ;
        RECT 95.420 14.250 95.790 14.260 ;
        RECT 99.265 14.170 100.290 14.430 ;
        RECT 100.745 14.260 101.770 14.520 ;
        RECT 105.245 14.430 105.615 14.440 ;
        RECT 100.745 14.250 101.115 14.260 ;
        RECT 104.590 14.170 105.615 14.430 ;
        RECT 106.080 14.260 107.105 14.520 ;
        RECT 110.580 14.430 110.950 14.440 ;
        RECT 106.080 14.250 106.450 14.260 ;
        RECT 109.925 14.170 110.950 14.430 ;
        RECT 111.405 14.260 112.430 14.520 ;
        RECT 115.905 14.430 116.275 14.440 ;
        RECT 111.405 14.250 111.775 14.260 ;
        RECT 115.250 14.170 116.275 14.430 ;
        RECT 116.740 14.260 117.765 14.520 ;
        RECT 121.240 14.430 121.610 14.440 ;
        RECT 116.740 14.250 117.110 14.260 ;
        RECT 120.585 14.170 121.610 14.430 ;
        RECT 41.285 14.160 41.655 14.170 ;
        RECT 46.620 14.160 46.990 14.170 ;
        RECT 51.945 14.160 52.315 14.170 ;
        RECT 57.280 14.160 57.650 14.170 ;
        RECT 62.605 14.160 62.975 14.170 ;
        RECT 67.940 14.160 68.310 14.170 ;
        RECT 73.265 14.160 73.635 14.170 ;
        RECT 78.600 14.160 78.970 14.170 ;
        RECT 83.925 14.160 84.295 14.170 ;
        RECT 89.260 14.160 89.630 14.170 ;
        RECT 94.585 14.160 94.955 14.170 ;
        RECT 99.920 14.160 100.290 14.170 ;
        RECT 105.245 14.160 105.615 14.170 ;
        RECT 110.580 14.160 110.950 14.170 ;
        RECT 115.905 14.160 116.275 14.170 ;
        RECT 121.240 14.160 121.610 14.170 ;
        RECT 28.410 12.475 28.690 12.845 ;
        RECT 36.785 12.495 37.155 12.505 ;
        RECT 42.120 12.495 42.490 12.505 ;
        RECT 47.445 12.495 47.815 12.505 ;
        RECT 52.780 12.495 53.150 12.505 ;
        RECT 58.105 12.495 58.475 12.505 ;
        RECT 63.440 12.495 63.810 12.505 ;
        RECT 68.765 12.495 69.135 12.505 ;
        RECT 74.100 12.495 74.470 12.505 ;
        RECT 79.425 12.495 79.795 12.505 ;
        RECT 84.760 12.495 85.130 12.505 ;
        RECT 90.085 12.495 90.455 12.505 ;
        RECT 95.420 12.495 95.790 12.505 ;
        RECT 100.745 12.495 101.115 12.505 ;
        RECT 106.080 12.495 106.450 12.505 ;
        RECT 111.405 12.495 111.775 12.505 ;
        RECT 116.740 12.495 117.110 12.505 ;
        RECT 28.035 11.180 28.315 11.550 ;
        RECT 27.325 11.000 27.505 11.045 ;
        RECT 25.375 10.540 25.655 10.910 ;
        RECT 28.085 8.730 28.265 11.180 ;
        RECT 10.530 3.080 10.790 8.595 ;
        RECT 11.745 8.075 13.345 8.365 ;
        RECT 12.430 2.525 12.690 8.075 ;
        RECT 16.040 7.630 17.645 7.920 ;
        RECT 16.110 7.070 16.565 7.630 ;
        RECT 28.045 7.625 28.305 8.730 ;
        RECT 15.455 6.615 16.565 7.070 ;
        RECT 15.455 3.610 15.910 6.615 ;
        RECT 28.465 4.435 28.645 12.475 ;
        RECT 36.785 12.235 37.810 12.495 ;
        RECT 41.285 12.400 41.655 12.410 ;
        RECT 36.785 12.225 37.155 12.235 ;
        RECT 40.630 12.140 41.655 12.400 ;
        RECT 42.120 12.235 43.145 12.495 ;
        RECT 46.620 12.400 46.990 12.410 ;
        RECT 42.120 12.225 42.490 12.235 ;
        RECT 45.965 12.140 46.330 12.400 ;
        RECT 46.575 12.140 46.990 12.400 ;
        RECT 47.445 12.235 48.470 12.495 ;
        RECT 51.945 12.400 52.315 12.410 ;
        RECT 47.445 12.225 47.815 12.235 ;
        RECT 51.290 12.140 52.315 12.400 ;
        RECT 52.780 12.235 53.805 12.495 ;
        RECT 57.280 12.400 57.650 12.410 ;
        RECT 52.780 12.225 53.150 12.235 ;
        RECT 56.625 12.140 56.990 12.400 ;
        RECT 57.235 12.140 57.650 12.400 ;
        RECT 58.105 12.235 59.130 12.495 ;
        RECT 62.605 12.400 62.975 12.410 ;
        RECT 58.105 12.225 58.475 12.235 ;
        RECT 61.950 12.140 62.975 12.400 ;
        RECT 63.440 12.235 64.465 12.495 ;
        RECT 67.940 12.400 68.310 12.410 ;
        RECT 63.440 12.225 63.810 12.235 ;
        RECT 67.285 12.140 67.650 12.400 ;
        RECT 67.895 12.140 68.310 12.400 ;
        RECT 68.765 12.235 69.790 12.495 ;
        RECT 73.265 12.400 73.635 12.410 ;
        RECT 68.765 12.225 69.135 12.235 ;
        RECT 72.610 12.140 73.635 12.400 ;
        RECT 74.100 12.235 75.125 12.495 ;
        RECT 78.600 12.400 78.970 12.410 ;
        RECT 74.100 12.225 74.470 12.235 ;
        RECT 77.945 12.140 78.310 12.400 ;
        RECT 78.555 12.140 78.970 12.400 ;
        RECT 79.425 12.235 80.450 12.495 ;
        RECT 83.925 12.400 84.295 12.410 ;
        RECT 79.425 12.225 79.795 12.235 ;
        RECT 83.270 12.140 84.295 12.400 ;
        RECT 84.760 12.235 85.785 12.495 ;
        RECT 89.260 12.400 89.630 12.410 ;
        RECT 84.760 12.225 85.130 12.235 ;
        RECT 88.605 12.140 88.970 12.400 ;
        RECT 89.215 12.140 89.630 12.400 ;
        RECT 90.085 12.235 91.110 12.495 ;
        RECT 94.585 12.400 94.955 12.410 ;
        RECT 90.085 12.225 90.455 12.235 ;
        RECT 93.930 12.140 94.955 12.400 ;
        RECT 95.420 12.235 96.445 12.495 ;
        RECT 99.920 12.400 100.290 12.410 ;
        RECT 95.420 12.225 95.790 12.235 ;
        RECT 99.265 12.140 99.630 12.400 ;
        RECT 99.875 12.140 100.290 12.400 ;
        RECT 100.745 12.235 101.770 12.495 ;
        RECT 105.245 12.400 105.615 12.410 ;
        RECT 100.745 12.225 101.115 12.235 ;
        RECT 104.590 12.140 105.615 12.400 ;
        RECT 106.080 12.235 107.105 12.495 ;
        RECT 110.580 12.400 110.950 12.410 ;
        RECT 106.080 12.225 106.450 12.235 ;
        RECT 109.925 12.140 110.290 12.400 ;
        RECT 110.535 12.140 110.950 12.400 ;
        RECT 111.405 12.235 112.430 12.495 ;
        RECT 115.905 12.400 116.275 12.410 ;
        RECT 111.405 12.225 111.775 12.235 ;
        RECT 115.250 12.140 116.275 12.400 ;
        RECT 116.740 12.235 117.765 12.495 ;
        RECT 121.240 12.400 121.610 12.410 ;
        RECT 116.740 12.225 117.110 12.235 ;
        RECT 120.585 12.140 120.950 12.400 ;
        RECT 121.195 12.140 121.610 12.400 ;
        RECT 41.285 12.130 41.655 12.140 ;
        RECT 34.005 11.845 34.400 11.850 ;
        RECT 33.390 11.565 35.160 11.845 ;
        RECT 38.715 11.565 39.110 11.845 ;
        RECT 39.330 11.570 39.740 11.850 ;
        RECT 40.020 11.565 40.485 11.845 ;
        RECT 44.050 11.565 44.445 11.845 ;
        RECT 44.665 11.570 45.075 11.850 ;
        RECT 45.355 11.565 45.820 11.845 ;
        RECT 46.010 11.505 46.255 12.140 ;
        RECT 46.620 12.130 46.990 12.140 ;
        RECT 51.945 12.130 52.315 12.140 ;
        RECT 49.375 11.565 49.770 11.845 ;
        RECT 49.990 11.570 50.400 11.850 ;
        RECT 50.680 11.565 51.145 11.845 ;
        RECT 54.710 11.565 55.105 11.845 ;
        RECT 55.325 11.570 55.735 11.850 ;
        RECT 56.015 11.565 56.480 11.845 ;
        RECT 56.670 11.505 56.915 12.140 ;
        RECT 57.280 12.130 57.650 12.140 ;
        RECT 62.605 12.130 62.975 12.140 ;
        RECT 60.035 11.565 60.430 11.845 ;
        RECT 60.650 11.570 61.060 11.850 ;
        RECT 61.340 11.565 61.805 11.845 ;
        RECT 65.370 11.565 65.765 11.845 ;
        RECT 65.985 11.570 66.395 11.850 ;
        RECT 66.675 11.565 67.140 11.845 ;
        RECT 67.330 11.505 67.575 12.140 ;
        RECT 67.940 12.130 68.310 12.140 ;
        RECT 73.265 12.130 73.635 12.140 ;
        RECT 70.695 11.565 71.090 11.845 ;
        RECT 71.310 11.570 71.720 11.850 ;
        RECT 72.000 11.565 72.465 11.845 ;
        RECT 76.030 11.565 76.425 11.845 ;
        RECT 76.645 11.570 77.055 11.850 ;
        RECT 77.335 11.565 77.800 11.845 ;
        RECT 77.990 11.505 78.235 12.140 ;
        RECT 78.600 12.130 78.970 12.140 ;
        RECT 83.925 12.130 84.295 12.140 ;
        RECT 81.355 11.565 81.750 11.845 ;
        RECT 81.970 11.570 82.380 11.850 ;
        RECT 82.660 11.565 83.125 11.845 ;
        RECT 86.690 11.565 87.085 11.845 ;
        RECT 87.305 11.570 87.715 11.850 ;
        RECT 87.995 11.565 88.460 11.845 ;
        RECT 88.650 11.505 88.895 12.140 ;
        RECT 89.260 12.130 89.630 12.140 ;
        RECT 94.585 12.130 94.955 12.140 ;
        RECT 92.015 11.565 92.410 11.845 ;
        RECT 92.630 11.570 93.040 11.850 ;
        RECT 93.320 11.565 93.785 11.845 ;
        RECT 97.350 11.565 97.745 11.845 ;
        RECT 97.965 11.570 98.375 11.850 ;
        RECT 98.655 11.565 99.120 11.845 ;
        RECT 99.310 11.505 99.555 12.140 ;
        RECT 99.920 12.130 100.290 12.140 ;
        RECT 105.245 12.130 105.615 12.140 ;
        RECT 102.675 11.565 103.070 11.845 ;
        RECT 103.290 11.570 103.700 11.850 ;
        RECT 103.980 11.565 104.445 11.845 ;
        RECT 108.010 11.565 108.405 11.845 ;
        RECT 108.625 11.570 109.035 11.850 ;
        RECT 109.315 11.565 109.780 11.845 ;
        RECT 109.970 11.505 110.215 12.140 ;
        RECT 110.580 12.130 110.950 12.140 ;
        RECT 115.905 12.130 116.275 12.140 ;
        RECT 113.335 11.565 113.730 11.845 ;
        RECT 113.950 11.570 114.360 11.850 ;
        RECT 114.640 11.565 115.105 11.845 ;
        RECT 118.670 11.565 119.065 11.845 ;
        RECT 119.285 11.570 119.695 11.850 ;
        RECT 119.975 11.565 120.440 11.845 ;
        RECT 120.630 11.505 120.875 12.140 ;
        RECT 121.240 12.130 121.610 12.140 ;
        RECT 124.610 11.845 125.005 11.850 ;
        RECT 123.995 11.565 125.765 11.845 ;
        RECT 46.010 11.260 46.930 11.505 ;
        RECT 56.670 11.260 57.590 11.505 ;
        RECT 67.330 11.260 68.250 11.505 ;
        RECT 77.990 11.260 78.910 11.505 ;
        RECT 88.650 11.260 89.570 11.505 ;
        RECT 99.310 11.260 100.230 11.505 ;
        RECT 109.970 11.260 110.890 11.505 ;
        RECT 120.630 11.260 121.550 11.505 ;
        RECT 36.785 11.195 37.155 11.205 ;
        RECT 42.120 11.195 42.490 11.205 ;
        RECT 36.785 10.935 37.860 11.195 ;
        RECT 42.120 10.935 43.195 11.195 ;
        RECT 36.785 10.925 37.155 10.935 ;
        RECT 42.120 10.925 42.490 10.935 ;
        RECT 46.685 10.575 46.930 11.260 ;
        RECT 47.445 11.195 47.815 11.205 ;
        RECT 52.780 11.195 53.150 11.205 ;
        RECT 47.445 10.935 48.520 11.195 ;
        RECT 52.780 10.935 53.855 11.195 ;
        RECT 47.445 10.925 47.815 10.935 ;
        RECT 52.780 10.925 53.150 10.935 ;
        RECT 57.345 10.575 57.590 11.260 ;
        RECT 58.105 11.195 58.475 11.205 ;
        RECT 63.440 11.195 63.810 11.205 ;
        RECT 58.105 10.935 59.180 11.195 ;
        RECT 63.440 10.935 64.515 11.195 ;
        RECT 58.105 10.925 58.475 10.935 ;
        RECT 63.440 10.925 63.810 10.935 ;
        RECT 68.005 10.575 68.250 11.260 ;
        RECT 68.765 11.195 69.135 11.205 ;
        RECT 74.100 11.195 74.470 11.205 ;
        RECT 68.765 10.935 69.840 11.195 ;
        RECT 74.100 10.935 75.175 11.195 ;
        RECT 68.765 10.925 69.135 10.935 ;
        RECT 74.100 10.925 74.470 10.935 ;
        RECT 78.665 10.575 78.910 11.260 ;
        RECT 79.425 11.195 79.795 11.205 ;
        RECT 84.760 11.195 85.130 11.205 ;
        RECT 79.425 10.935 80.500 11.195 ;
        RECT 84.760 10.935 85.835 11.195 ;
        RECT 79.425 10.925 79.795 10.935 ;
        RECT 84.760 10.925 85.130 10.935 ;
        RECT 89.325 10.575 89.570 11.260 ;
        RECT 90.085 11.195 90.455 11.205 ;
        RECT 95.420 11.195 95.790 11.205 ;
        RECT 90.085 10.935 91.160 11.195 ;
        RECT 95.420 10.935 96.495 11.195 ;
        RECT 90.085 10.925 90.455 10.935 ;
        RECT 95.420 10.925 95.790 10.935 ;
        RECT 99.985 10.575 100.230 11.260 ;
        RECT 100.745 11.195 101.115 11.205 ;
        RECT 106.080 11.195 106.450 11.205 ;
        RECT 100.745 10.935 101.820 11.195 ;
        RECT 106.080 10.935 107.155 11.195 ;
        RECT 100.745 10.925 101.115 10.935 ;
        RECT 106.080 10.925 106.450 10.935 ;
        RECT 110.645 10.575 110.890 11.260 ;
        RECT 111.405 11.195 111.775 11.205 ;
        RECT 116.740 11.195 117.110 11.205 ;
        RECT 111.405 10.935 112.480 11.195 ;
        RECT 116.740 10.935 117.815 11.195 ;
        RECT 111.405 10.925 111.775 10.935 ;
        RECT 116.740 10.925 117.110 10.935 ;
        RECT 121.305 10.575 121.550 11.260 ;
        RECT 41.290 10.565 41.660 10.575 ;
        RECT 40.630 10.305 41.660 10.565 ;
        RECT 41.290 10.295 41.660 10.305 ;
        RECT 45.940 10.290 46.360 10.570 ;
        RECT 46.625 10.295 46.995 10.575 ;
        RECT 51.950 10.565 52.320 10.575 ;
        RECT 51.290 10.305 52.320 10.565 ;
        RECT 51.950 10.295 52.320 10.305 ;
        RECT 56.600 10.290 57.020 10.570 ;
        RECT 57.285 10.295 57.655 10.575 ;
        RECT 62.610 10.565 62.980 10.575 ;
        RECT 61.950 10.305 62.980 10.565 ;
        RECT 62.610 10.295 62.980 10.305 ;
        RECT 67.260 10.290 67.680 10.570 ;
        RECT 67.945 10.295 68.315 10.575 ;
        RECT 73.270 10.565 73.640 10.575 ;
        RECT 72.610 10.305 73.640 10.565 ;
        RECT 73.270 10.295 73.640 10.305 ;
        RECT 77.920 10.290 78.340 10.570 ;
        RECT 78.605 10.295 78.975 10.575 ;
        RECT 83.930 10.565 84.300 10.575 ;
        RECT 83.270 10.305 84.300 10.565 ;
        RECT 83.930 10.295 84.300 10.305 ;
        RECT 88.580 10.290 89.000 10.570 ;
        RECT 89.265 10.295 89.635 10.575 ;
        RECT 94.590 10.565 94.960 10.575 ;
        RECT 93.930 10.305 94.960 10.565 ;
        RECT 94.590 10.295 94.960 10.305 ;
        RECT 99.240 10.290 99.660 10.570 ;
        RECT 99.925 10.295 100.295 10.575 ;
        RECT 105.250 10.565 105.620 10.575 ;
        RECT 104.590 10.305 105.620 10.565 ;
        RECT 105.250 10.295 105.620 10.305 ;
        RECT 109.900 10.290 110.320 10.570 ;
        RECT 110.585 10.295 110.955 10.575 ;
        RECT 115.910 10.565 116.280 10.575 ;
        RECT 115.250 10.305 116.280 10.565 ;
        RECT 115.910 10.295 116.280 10.305 ;
        RECT 120.560 10.290 120.980 10.570 ;
        RECT 121.245 10.295 121.615 10.575 ;
        RECT 32.625 7.205 34.390 7.485 ;
        RECT 37.950 7.205 39.715 7.485 ;
        RECT 43.285 7.205 45.050 7.485 ;
        RECT 48.610 7.205 50.375 7.485 ;
        RECT 53.945 7.205 55.710 7.485 ;
        RECT 59.270 7.205 61.035 7.485 ;
        RECT 64.605 7.205 66.370 7.485 ;
        RECT 69.930 7.205 71.695 7.485 ;
        RECT 75.265 7.205 77.030 7.485 ;
        RECT 80.590 7.205 82.355 7.485 ;
        RECT 85.925 7.205 87.690 7.485 ;
        RECT 91.250 7.205 93.015 7.485 ;
        RECT 96.585 7.205 98.350 7.485 ;
        RECT 101.910 7.205 103.675 7.485 ;
        RECT 107.245 7.205 109.010 7.485 ;
        RECT 112.570 7.205 114.335 7.485 ;
        RECT 117.905 7.205 119.670 7.485 ;
        RECT 123.230 7.205 124.995 7.485 ;
        RECT 28.465 4.280 28.655 4.435 ;
        RECT 34.005 4.310 34.400 4.315 ;
        RECT 38.900 4.310 40.145 4.315 ;
        RECT 44.275 4.310 45.460 4.315 ;
        RECT 49.560 4.310 50.805 4.315 ;
        RECT 54.935 4.310 56.120 4.315 ;
        RECT 60.220 4.310 61.465 4.315 ;
        RECT 65.595 4.310 66.780 4.315 ;
        RECT 70.880 4.310 72.125 4.315 ;
        RECT 76.255 4.310 77.440 4.315 ;
        RECT 81.540 4.310 82.785 4.315 ;
        RECT 86.915 4.310 88.100 4.315 ;
        RECT 92.200 4.310 93.445 4.315 ;
        RECT 97.575 4.310 98.760 4.315 ;
        RECT 102.860 4.310 104.105 4.315 ;
        RECT 108.235 4.310 109.420 4.315 ;
        RECT 113.520 4.310 114.765 4.315 ;
        RECT 118.895 4.310 120.080 4.315 ;
        RECT 124.610 4.310 125.005 4.315 ;
        RECT 28.475 4.010 28.655 4.280 ;
        RECT 33.390 4.030 35.160 4.310 ;
        RECT 38.715 4.035 40.485 4.310 ;
        RECT 38.715 4.030 39.110 4.035 ;
        RECT 40.120 4.030 40.485 4.035 ;
        RECT 44.050 4.035 45.820 4.310 ;
        RECT 44.050 4.030 44.445 4.035 ;
        RECT 45.455 4.030 45.820 4.035 ;
        RECT 49.375 4.035 51.145 4.310 ;
        RECT 49.375 4.030 49.770 4.035 ;
        RECT 50.780 4.030 51.145 4.035 ;
        RECT 54.710 4.035 56.480 4.310 ;
        RECT 54.710 4.030 55.105 4.035 ;
        RECT 56.115 4.030 56.480 4.035 ;
        RECT 60.035 4.035 61.805 4.310 ;
        RECT 60.035 4.030 60.430 4.035 ;
        RECT 61.440 4.030 61.805 4.035 ;
        RECT 65.370 4.035 67.140 4.310 ;
        RECT 65.370 4.030 65.765 4.035 ;
        RECT 66.775 4.030 67.140 4.035 ;
        RECT 70.695 4.035 72.465 4.310 ;
        RECT 70.695 4.030 71.090 4.035 ;
        RECT 72.100 4.030 72.465 4.035 ;
        RECT 76.030 4.035 77.800 4.310 ;
        RECT 76.030 4.030 76.425 4.035 ;
        RECT 77.435 4.030 77.800 4.035 ;
        RECT 81.355 4.035 83.125 4.310 ;
        RECT 81.355 4.030 81.750 4.035 ;
        RECT 82.760 4.030 83.125 4.035 ;
        RECT 86.690 4.035 88.460 4.310 ;
        RECT 86.690 4.030 87.085 4.035 ;
        RECT 88.095 4.030 88.460 4.035 ;
        RECT 92.015 4.035 93.785 4.310 ;
        RECT 92.015 4.030 92.410 4.035 ;
        RECT 93.420 4.030 93.785 4.035 ;
        RECT 97.350 4.035 99.120 4.310 ;
        RECT 97.350 4.030 97.745 4.035 ;
        RECT 98.755 4.030 99.120 4.035 ;
        RECT 102.675 4.035 104.445 4.310 ;
        RECT 102.675 4.030 103.070 4.035 ;
        RECT 104.080 4.030 104.445 4.035 ;
        RECT 108.010 4.035 109.780 4.310 ;
        RECT 108.010 4.030 108.405 4.035 ;
        RECT 109.415 4.030 109.780 4.035 ;
        RECT 113.335 4.035 115.105 4.310 ;
        RECT 113.335 4.030 113.730 4.035 ;
        RECT 114.740 4.030 115.105 4.035 ;
        RECT 118.670 4.035 120.440 4.310 ;
        RECT 118.670 4.030 119.065 4.035 ;
        RECT 120.075 4.030 120.440 4.035 ;
        RECT 123.995 4.030 125.765 4.310 ;
        RECT 14.605 3.320 15.985 3.610 ;
        RECT 28.435 2.905 28.695 4.010 ;
        RECT 28.475 2.860 28.655 2.905 ;
      LAYER met3 ;
        RECT 53.470 80.860 53.770 81.275 ;
        RECT 42.810 80.100 43.110 80.515 ;
        RECT 53.455 80.510 53.785 80.860 ;
        RECT 42.795 79.750 43.125 80.100 ;
        RECT 38.760 69.835 39.060 70.230 ;
        RECT 24.575 68.825 24.925 68.840 ;
        RECT 29.710 68.825 30.960 68.835 ;
        RECT 24.575 68.525 30.975 68.825 ;
        RECT 36.810 68.795 37.140 69.600 ;
        RECT 38.750 69.455 39.070 69.835 ;
        RECT 42.810 69.820 43.110 79.750 ;
        RECT 43.440 79.710 43.740 80.125 ;
        RECT 43.425 79.360 43.755 79.710 ;
        RECT 42.145 69.520 43.110 69.820 ;
        RECT 24.575 68.510 24.925 68.525 ;
        RECT 29.710 68.515 30.960 68.525 ;
        RECT 36.810 68.485 37.130 68.795 ;
        RECT 28.000 68.180 28.350 68.195 ;
        RECT 29.710 68.180 30.960 68.190 ;
        RECT 27.975 67.880 30.975 68.180 ;
        RECT 28.000 67.865 28.350 67.880 ;
        RECT 29.710 67.870 30.960 67.880 ;
        RECT 36.820 67.670 37.120 67.970 ;
        RECT 38.760 67.800 39.060 69.455 ;
        RECT 42.145 68.795 42.475 69.520 ;
        RECT 43.440 68.495 43.740 79.360 ;
        RECT 44.085 73.385 44.405 73.765 ;
        RECT 24.200 67.535 24.550 67.550 ;
        RECT 29.710 67.535 30.960 67.545 ;
        RECT 24.200 67.235 30.975 67.535 ;
        RECT 24.200 67.220 24.550 67.235 ;
        RECT 29.710 67.225 30.960 67.235 ;
        RECT 36.805 66.935 37.135 67.670 ;
        RECT 37.970 67.450 38.300 67.800 ;
        RECT 38.745 67.450 39.075 67.800 ;
        RECT 39.380 67.450 39.710 67.800 ;
        RECT 41.305 67.535 41.635 68.270 ;
        RECT 42.140 68.195 43.740 68.495 ;
        RECT 28.380 66.890 28.730 66.905 ;
        RECT 29.710 66.890 30.960 66.900 ;
        RECT 28.355 66.590 30.975 66.890 ;
        RECT 28.380 66.575 28.730 66.590 ;
        RECT 29.710 66.580 30.960 66.590 ;
        RECT 37.985 66.300 38.285 67.450 ;
        RECT 37.975 65.920 38.295 66.300 ;
        RECT 27.995 65.560 28.345 65.575 ;
        RECT 27.995 65.555 28.760 65.560 ;
        RECT 29.710 65.555 30.960 65.565 ;
        RECT 27.965 65.255 30.975 65.555 ;
        RECT 27.995 65.245 28.345 65.255 ;
        RECT 29.710 65.245 30.960 65.255 ;
        RECT 27.240 64.910 27.590 64.925 ;
        RECT 36.805 64.920 37.135 65.670 ;
        RECT 29.710 64.910 30.960 64.920 ;
        RECT 27.200 64.610 30.975 64.910 ;
        RECT 39.395 64.630 39.695 67.450 ;
        RECT 41.305 66.485 41.635 67.235 ;
        RECT 42.140 66.935 42.470 68.195 ;
        RECT 44.095 67.800 44.395 73.385 ;
        RECT 49.420 69.835 49.720 70.230 ;
        RECT 47.470 69.145 47.800 69.600 ;
        RECT 49.410 69.455 49.730 69.835 ;
        RECT 53.470 69.820 53.770 80.510 ;
        RECT 54.100 80.470 54.400 80.885 ;
        RECT 54.085 80.120 54.415 80.470 ;
        RECT 52.805 69.520 53.770 69.820 ;
        RECT 45.790 68.845 47.800 69.145 ;
        RECT 43.305 67.450 43.635 67.800 ;
        RECT 44.080 67.450 44.410 67.800 ;
        RECT 44.715 67.450 45.045 67.800 ;
        RECT 45.790 67.575 46.090 68.845 ;
        RECT 47.470 68.795 47.800 68.845 ;
        RECT 48.100 68.485 48.420 68.865 ;
        RECT 48.100 68.390 48.410 68.485 ;
        RECT 43.320 66.300 43.620 67.450 ;
        RECT 43.310 65.920 43.630 66.300 ;
        RECT 27.240 64.595 27.590 64.610 ;
        RECT 29.710 64.600 30.960 64.610 ;
        RECT 28.380 64.265 28.730 64.280 ;
        RECT 29.710 64.265 30.960 64.275 ;
        RECT 28.350 63.965 30.975 64.265 ;
        RECT 28.380 63.950 28.730 63.965 ;
        RECT 29.710 63.955 30.960 63.965 ;
        RECT 27.620 63.620 27.970 63.635 ;
        RECT 29.710 63.620 30.960 63.630 ;
        RECT 36.805 63.620 37.135 64.370 ;
        RECT 38.750 64.275 39.080 64.625 ;
        RECT 39.380 64.280 39.710 64.630 ;
        RECT 27.605 63.320 30.975 63.620 ;
        RECT 27.620 63.305 27.970 63.320 ;
        RECT 29.710 63.310 30.960 63.320 ;
        RECT 27.235 61.290 27.585 61.305 ;
        RECT 29.710 61.290 30.960 61.300 ;
        RECT 27.220 60.990 30.975 61.290 ;
        RECT 27.235 60.975 27.585 60.990 ;
        RECT 29.710 60.980 30.960 60.990 ;
        RECT 36.810 60.885 37.140 61.635 ;
        RECT 28.380 60.645 28.730 60.660 ;
        RECT 29.710 60.645 30.960 60.655 ;
        RECT 28.335 60.345 30.975 60.645 ;
        RECT 28.380 60.330 28.730 60.345 ;
        RECT 29.710 60.335 30.960 60.345 ;
        RECT 38.765 60.265 39.065 64.275 ;
        RECT 39.395 60.265 39.695 64.280 ;
        RECT 40.035 64.275 40.365 64.625 ;
        RECT 41.305 64.435 41.635 65.195 ;
        RECT 42.140 64.920 42.470 65.670 ;
        RECT 44.730 64.630 45.030 67.450 ;
        RECT 45.780 67.195 46.100 67.575 ;
        RECT 46.640 67.535 46.970 68.270 ;
        RECT 47.465 68.090 48.410 68.390 ;
        RECT 46.640 66.485 46.970 67.235 ;
        RECT 47.465 66.935 47.795 68.090 ;
        RECT 49.420 67.800 49.720 69.455 ;
        RECT 52.805 68.795 53.135 69.520 ;
        RECT 54.100 68.495 54.400 80.120 ;
        RECT 64.130 79.720 64.430 80.135 ;
        RECT 64.760 80.090 65.060 80.505 ;
        RECT 85.450 80.100 85.750 80.515 ;
        RECT 96.110 80.480 96.410 80.895 ;
        RECT 96.725 80.515 97.055 80.865 ;
        RECT 96.095 80.130 96.425 80.480 ;
        RECT 64.745 79.740 65.075 80.090 ;
        RECT 85.435 79.750 85.765 80.100 ;
        RECT 64.115 79.370 64.445 79.720 ;
        RECT 54.745 73.385 55.065 73.765 ;
        RECT 48.630 67.450 48.960 67.800 ;
        RECT 49.405 67.450 49.735 67.800 ;
        RECT 50.040 67.450 50.370 67.800 ;
        RECT 51.965 67.535 52.295 68.270 ;
        RECT 52.800 68.195 54.400 68.495 ;
        RECT 48.645 66.300 48.945 67.450 ;
        RECT 48.635 65.920 48.955 66.300 ;
        RECT 27.620 60.000 27.970 60.015 ;
        RECT 29.710 60.000 30.960 60.010 ;
        RECT 27.590 59.700 30.975 60.000 ;
        RECT 27.620 59.685 27.970 59.700 ;
        RECT 29.710 59.690 30.960 59.700 ;
        RECT 28.000 59.355 28.350 59.370 ;
        RECT 29.710 59.355 30.960 59.365 ;
        RECT 27.975 59.055 30.975 59.355 ;
        RECT 36.805 59.350 37.135 60.105 ;
        RECT 38.120 59.915 38.450 60.265 ;
        RECT 38.750 59.915 39.080 60.265 ;
        RECT 39.380 59.915 39.710 60.265 ;
        RECT 28.000 59.040 28.350 59.055 ;
        RECT 29.710 59.045 30.960 59.055 ;
        RECT 28.375 58.025 28.725 58.040 ;
        RECT 28.375 58.020 29.140 58.025 ;
        RECT 29.710 58.020 30.960 58.030 ;
        RECT 28.355 57.720 30.975 58.020 ;
        RECT 28.375 57.710 28.725 57.720 ;
        RECT 29.710 57.710 30.960 57.720 ;
        RECT 26.480 57.375 26.830 57.390 ;
        RECT 36.805 57.385 37.135 58.135 ;
        RECT 29.710 57.375 30.960 57.385 ;
        RECT 26.470 57.075 30.975 57.375 ;
        RECT 26.480 57.060 26.830 57.075 ;
        RECT 29.710 57.065 30.960 57.075 ;
        RECT 28.000 56.730 28.350 56.745 ;
        RECT 29.710 56.730 30.960 56.740 ;
        RECT 27.985 56.430 30.975 56.730 ;
        RECT 28.000 56.415 28.350 56.430 ;
        RECT 29.710 56.420 30.960 56.430 ;
        RECT 26.860 56.085 27.210 56.100 ;
        RECT 29.710 56.085 30.960 56.095 ;
        RECT 36.805 56.085 37.135 56.835 ;
        RECT 26.835 55.785 30.975 56.085 ;
        RECT 26.860 55.770 27.210 55.785 ;
        RECT 29.710 55.775 30.960 55.785 ;
        RECT 26.475 53.755 26.825 53.770 ;
        RECT 29.710 53.755 30.960 53.765 ;
        RECT 26.435 53.455 30.975 53.755 ;
        RECT 26.475 53.440 26.825 53.455 ;
        RECT 29.710 53.445 30.960 53.455 ;
        RECT 36.810 53.350 37.140 54.100 ;
        RECT 28.000 53.110 28.350 53.125 ;
        RECT 29.710 53.110 30.960 53.120 ;
        RECT 27.970 52.810 30.975 53.110 ;
        RECT 37.450 52.960 37.780 53.310 ;
        RECT 38.135 53.145 38.435 59.915 ;
        RECT 38.765 57.090 39.065 59.915 ;
        RECT 40.050 57.505 40.350 64.275 ;
        RECT 41.310 62.990 41.640 63.740 ;
        RECT 42.140 63.620 42.470 64.370 ;
        RECT 44.085 64.275 44.415 64.625 ;
        RECT 44.715 64.280 45.045 64.630 ;
        RECT 41.305 60.235 41.635 60.985 ;
        RECT 42.145 60.885 42.475 61.635 ;
        RECT 44.100 60.265 44.400 64.275 ;
        RECT 44.730 60.265 45.030 64.280 ;
        RECT 45.370 64.275 45.700 64.625 ;
        RECT 46.640 64.435 46.970 65.195 ;
        RECT 47.465 64.920 47.795 65.670 ;
        RECT 50.055 64.630 50.355 67.450 ;
        RECT 51.965 66.485 52.295 67.235 ;
        RECT 52.800 66.935 53.130 68.195 ;
        RECT 54.755 67.800 55.055 73.385 ;
        RECT 60.080 69.835 60.380 70.230 ;
        RECT 58.130 68.795 58.460 69.600 ;
        RECT 60.070 69.455 60.390 69.835 ;
        RECT 64.130 69.820 64.430 79.370 ;
        RECT 63.465 69.520 64.430 69.820 ;
        RECT 58.130 68.485 58.450 68.795 ;
        RECT 54.740 67.450 55.070 67.800 ;
        RECT 55.375 67.450 55.705 67.800 ;
        RECT 57.300 67.535 57.630 68.270 ;
        RECT 58.140 67.670 58.440 67.970 ;
        RECT 60.080 67.800 60.380 69.455 ;
        RECT 63.465 68.795 63.795 69.520 ;
        RECT 64.760 68.495 65.060 79.740 ;
        RECT 65.405 73.385 65.725 73.765 ;
        RECT 41.305 58.950 41.635 59.700 ;
        RECT 42.140 59.350 42.470 60.105 ;
        RECT 43.455 59.915 43.785 60.265 ;
        RECT 44.085 59.915 44.415 60.265 ;
        RECT 44.715 59.915 45.045 60.265 ;
        RECT 40.050 57.090 40.365 57.505 ;
        RECT 38.750 56.740 39.080 57.090 ;
        RECT 40.050 56.740 40.380 57.090 ;
        RECT 41.305 56.900 41.635 57.660 ;
        RECT 42.140 57.385 42.470 58.135 ;
        RECT 28.000 52.795 28.350 52.810 ;
        RECT 29.710 52.800 30.960 52.810 ;
        RECT 26.860 52.465 27.210 52.480 ;
        RECT 29.710 52.465 30.960 52.475 ;
        RECT 26.845 52.165 30.975 52.465 ;
        RECT 26.860 52.150 27.210 52.165 ;
        RECT 29.710 52.155 30.960 52.165 ;
        RECT 28.380 51.820 28.730 51.835 ;
        RECT 29.710 51.820 30.960 51.830 ;
        RECT 28.350 51.520 30.975 51.820 ;
        RECT 36.805 51.815 37.135 52.570 ;
        RECT 28.380 51.505 28.730 51.520 ;
        RECT 29.710 51.510 30.960 51.520 ;
        RECT 27.995 50.490 28.345 50.505 ;
        RECT 27.995 50.485 28.760 50.490 ;
        RECT 29.710 50.485 30.960 50.495 ;
        RECT 27.970 50.185 30.975 50.485 ;
        RECT 27.995 50.175 28.345 50.185 ;
        RECT 29.710 50.175 30.960 50.185 ;
        RECT 27.620 49.840 27.970 49.855 ;
        RECT 36.805 49.850 37.135 50.600 ;
        RECT 29.710 49.840 30.960 49.850 ;
        RECT 27.585 49.540 30.975 49.840 ;
        RECT 27.620 49.525 27.970 49.540 ;
        RECT 29.710 49.530 30.960 49.540 ;
        RECT 28.380 49.195 28.730 49.210 ;
        RECT 29.710 49.195 30.960 49.205 ;
        RECT 28.350 48.895 30.975 49.195 ;
        RECT 28.380 48.880 28.730 48.895 ;
        RECT 29.710 48.885 30.960 48.895 ;
        RECT 27.240 48.550 27.590 48.565 ;
        RECT 29.710 48.550 30.960 48.560 ;
        RECT 36.805 48.550 37.135 49.300 ;
        RECT 27.230 48.250 30.975 48.550 ;
        RECT 27.240 48.235 27.590 48.250 ;
        RECT 29.710 48.240 30.960 48.250 ;
        RECT 27.615 46.220 27.965 46.235 ;
        RECT 29.710 46.220 30.960 46.230 ;
        RECT 27.585 45.920 30.975 46.220 ;
        RECT 27.615 45.905 27.965 45.920 ;
        RECT 29.710 45.910 30.960 45.920 ;
        RECT 36.810 45.815 37.140 46.565 ;
        RECT 28.380 45.575 28.730 45.590 ;
        RECT 29.710 45.575 30.960 45.585 ;
        RECT 28.350 45.275 30.975 45.575 ;
        RECT 28.380 45.260 28.730 45.275 ;
        RECT 29.710 45.265 30.960 45.275 ;
        RECT 27.240 44.930 27.590 44.945 ;
        RECT 29.710 44.930 30.960 44.940 ;
        RECT 27.215 44.630 30.975 44.930 ;
        RECT 27.240 44.615 27.590 44.630 ;
        RECT 29.710 44.620 30.960 44.630 ;
        RECT 28.000 44.285 28.350 44.300 ;
        RECT 29.710 44.285 30.960 44.295 ;
        RECT 27.970 43.985 30.975 44.285 ;
        RECT 36.805 44.280 37.135 45.035 ;
        RECT 28.000 43.970 28.350 43.985 ;
        RECT 29.710 43.975 30.960 43.985 ;
        RECT 28.375 42.955 28.725 42.970 ;
        RECT 28.375 42.950 29.140 42.955 ;
        RECT 29.710 42.950 30.960 42.960 ;
        RECT 28.340 42.650 30.975 42.950 ;
        RECT 28.375 42.640 28.725 42.650 ;
        RECT 29.710 42.640 30.960 42.650 ;
        RECT 26.100 42.305 26.450 42.320 ;
        RECT 36.805 42.315 37.135 43.065 ;
        RECT 29.710 42.305 30.960 42.315 ;
        RECT 26.060 42.005 30.975 42.305 ;
        RECT 26.100 41.990 26.450 42.005 ;
        RECT 29.710 41.995 30.960 42.005 ;
        RECT 28.000 41.660 28.350 41.675 ;
        RECT 29.710 41.660 30.960 41.670 ;
        RECT 27.970 41.360 30.975 41.660 ;
        RECT 28.000 41.345 28.350 41.360 ;
        RECT 29.710 41.350 30.960 41.360 ;
        RECT 25.720 41.015 26.070 41.030 ;
        RECT 29.710 41.015 30.960 41.025 ;
        RECT 36.805 41.015 37.135 41.765 ;
        RECT 25.710 40.715 30.975 41.015 ;
        RECT 25.720 40.700 26.070 40.715 ;
        RECT 29.710 40.705 30.960 40.715 ;
        RECT 26.095 38.685 26.445 38.700 ;
        RECT 29.710 38.685 30.960 38.695 ;
        RECT 26.065 38.385 30.975 38.685 ;
        RECT 26.095 38.370 26.445 38.385 ;
        RECT 29.710 38.375 30.960 38.385 ;
        RECT 36.810 38.280 37.140 39.030 ;
        RECT 28.000 38.040 28.350 38.055 ;
        RECT 29.710 38.040 30.960 38.050 ;
        RECT 27.970 37.740 30.975 38.040 ;
        RECT 28.000 37.725 28.350 37.740 ;
        RECT 29.710 37.730 30.960 37.740 ;
        RECT 37.465 37.660 37.765 52.960 ;
        RECT 38.135 52.730 38.450 53.145 ;
        RECT 38.135 52.380 38.465 52.730 ;
        RECT 39.380 52.380 39.710 52.730 ;
        RECT 38.135 45.195 38.435 52.380 ;
        RECT 39.395 49.560 39.695 52.380 ;
        RECT 38.750 49.205 39.080 49.555 ;
        RECT 39.380 49.210 39.710 49.560 ;
        RECT 40.050 49.555 40.350 56.740 ;
        RECT 40.665 56.235 40.995 56.585 ;
        RECT 38.765 45.195 39.065 49.205 ;
        RECT 39.395 45.195 39.695 49.210 ;
        RECT 40.035 49.205 40.365 49.555 ;
        RECT 38.120 44.845 38.450 45.195 ;
        RECT 38.750 44.845 39.080 45.195 ;
        RECT 39.380 44.845 39.710 45.195 ;
        RECT 38.765 42.020 39.065 44.845 ;
        RECT 38.750 41.670 39.080 42.020 ;
        RECT 39.405 41.675 39.735 42.025 ;
        RECT 40.680 42.020 40.980 56.235 ;
        RECT 41.310 55.455 41.640 56.205 ;
        RECT 42.140 56.085 42.470 56.835 ;
        RECT 41.305 52.700 41.635 53.450 ;
        RECT 42.145 53.350 42.475 54.100 ;
        RECT 42.785 52.960 43.115 53.310 ;
        RECT 43.470 53.145 43.770 59.915 ;
        RECT 44.100 57.090 44.400 59.915 ;
        RECT 45.385 57.505 45.685 64.275 ;
        RECT 46.645 62.990 46.975 63.740 ;
        RECT 47.465 63.620 47.795 64.370 ;
        RECT 49.410 64.275 49.740 64.625 ;
        RECT 50.040 64.280 50.370 64.630 ;
        RECT 46.640 60.235 46.970 60.985 ;
        RECT 47.470 60.885 47.800 61.635 ;
        RECT 49.425 60.265 49.725 64.275 ;
        RECT 50.055 60.265 50.355 64.280 ;
        RECT 50.695 64.275 51.025 64.625 ;
        RECT 51.965 64.435 52.295 65.195 ;
        RECT 52.800 64.920 53.130 65.670 ;
        RECT 55.390 64.630 55.690 67.450 ;
        RECT 57.300 66.485 57.630 67.235 ;
        RECT 58.125 66.935 58.455 67.670 ;
        RECT 59.290 67.450 59.620 67.800 ;
        RECT 60.065 67.450 60.395 67.800 ;
        RECT 60.700 67.450 61.030 67.800 ;
        RECT 62.625 67.535 62.955 68.270 ;
        RECT 63.460 68.195 65.060 68.495 ;
        RECT 59.305 66.300 59.605 67.450 ;
        RECT 59.295 65.920 59.615 66.300 ;
        RECT 46.640 58.950 46.970 59.700 ;
        RECT 47.465 59.350 47.795 60.105 ;
        RECT 48.780 59.915 49.110 60.265 ;
        RECT 49.410 59.915 49.740 60.265 ;
        RECT 50.040 59.915 50.370 60.265 ;
        RECT 45.385 57.090 45.700 57.505 ;
        RECT 44.085 56.740 44.415 57.090 ;
        RECT 45.385 56.740 45.715 57.090 ;
        RECT 46.640 56.900 46.970 57.660 ;
        RECT 47.465 57.385 47.795 58.135 ;
        RECT 41.305 51.415 41.635 52.165 ;
        RECT 42.140 51.815 42.470 52.570 ;
        RECT 41.305 49.365 41.635 50.125 ;
        RECT 42.140 49.850 42.470 50.600 ;
        RECT 41.310 47.920 41.640 48.670 ;
        RECT 42.140 48.550 42.470 49.300 ;
        RECT 41.305 45.165 41.635 45.915 ;
        RECT 42.145 45.815 42.475 46.565 ;
        RECT 41.305 43.880 41.635 44.630 ;
        RECT 42.140 44.280 42.470 45.035 ;
        RECT 25.720 37.395 26.070 37.410 ;
        RECT 29.710 37.395 30.960 37.405 ;
        RECT 25.695 37.095 30.975 37.395 ;
        RECT 25.720 37.080 26.070 37.095 ;
        RECT 29.710 37.085 30.960 37.095 ;
        RECT 28.380 36.750 28.730 36.765 ;
        RECT 29.710 36.750 30.960 36.760 ;
        RECT 28.325 36.450 30.975 36.750 ;
        RECT 36.805 36.745 37.135 37.500 ;
        RECT 37.450 37.310 37.780 37.660 ;
        RECT 28.380 36.435 28.730 36.450 ;
        RECT 29.710 36.440 30.960 36.450 ;
        RECT 27.995 35.420 28.345 35.435 ;
        RECT 27.995 35.415 28.760 35.420 ;
        RECT 29.710 35.415 30.960 35.425 ;
        RECT 27.965 35.115 30.975 35.415 ;
        RECT 27.995 35.105 28.345 35.115 ;
        RECT 29.710 35.105 30.960 35.115 ;
        RECT 27.240 34.770 27.590 34.785 ;
        RECT 36.805 34.780 37.135 35.530 ;
        RECT 29.710 34.770 30.960 34.780 ;
        RECT 27.205 34.470 30.975 34.770 ;
        RECT 27.240 34.455 27.590 34.470 ;
        RECT 29.710 34.460 30.960 34.470 ;
        RECT 28.380 34.125 28.730 34.140 ;
        RECT 29.710 34.125 30.960 34.135 ;
        RECT 28.355 33.825 30.975 34.125 ;
        RECT 28.380 33.810 28.730 33.825 ;
        RECT 29.710 33.815 30.960 33.825 ;
        RECT 27.620 33.480 27.970 33.495 ;
        RECT 29.710 33.480 30.960 33.490 ;
        RECT 36.805 33.480 37.135 34.230 ;
        RECT 27.585 33.180 30.975 33.480 ;
        RECT 27.620 33.165 27.970 33.180 ;
        RECT 29.710 33.170 30.960 33.180 ;
        RECT 27.235 31.150 27.585 31.165 ;
        RECT 29.710 31.150 30.960 31.160 ;
        RECT 27.220 30.850 30.975 31.150 ;
        RECT 27.235 30.835 27.585 30.850 ;
        RECT 29.710 30.840 30.960 30.850 ;
        RECT 36.810 30.745 37.140 31.495 ;
        RECT 28.380 30.505 28.730 30.520 ;
        RECT 29.710 30.505 30.960 30.515 ;
        RECT 28.355 30.205 30.975 30.505 ;
        RECT 28.380 30.190 28.730 30.205 ;
        RECT 29.710 30.195 30.960 30.205 ;
        RECT 27.620 29.860 27.970 29.875 ;
        RECT 29.710 29.860 30.960 29.870 ;
        RECT 27.580 29.560 30.975 29.860 ;
        RECT 27.620 29.545 27.970 29.560 ;
        RECT 29.710 29.550 30.960 29.560 ;
        RECT 28.000 29.215 28.350 29.230 ;
        RECT 29.710 29.215 30.960 29.225 ;
        RECT 27.955 28.915 30.975 29.215 ;
        RECT 36.805 29.210 37.135 29.965 ;
        RECT 28.000 28.900 28.350 28.915 ;
        RECT 29.710 28.905 30.960 28.915 ;
        RECT 28.375 27.885 28.725 27.900 ;
        RECT 28.375 27.880 29.140 27.885 ;
        RECT 29.710 27.880 30.960 27.890 ;
        RECT 28.355 27.580 30.975 27.880 ;
        RECT 28.375 27.570 28.725 27.580 ;
        RECT 29.710 27.570 30.960 27.580 ;
        RECT 26.860 27.235 27.210 27.250 ;
        RECT 36.805 27.245 37.135 27.995 ;
        RECT 29.710 27.235 30.960 27.245 ;
        RECT 26.850 26.935 30.975 27.235 ;
        RECT 26.860 26.920 27.210 26.935 ;
        RECT 29.710 26.925 30.960 26.935 ;
        RECT 28.000 26.590 28.350 26.605 ;
        RECT 29.710 26.590 30.960 26.600 ;
        RECT 27.970 26.290 30.975 26.590 ;
        RECT 28.000 26.275 28.350 26.290 ;
        RECT 29.710 26.280 30.960 26.290 ;
        RECT 26.480 25.945 26.830 25.960 ;
        RECT 29.710 25.945 30.960 25.955 ;
        RECT 36.805 25.945 37.135 26.695 ;
        RECT 26.465 25.645 30.975 25.945 ;
        RECT 26.480 25.630 26.830 25.645 ;
        RECT 29.710 25.635 30.960 25.645 ;
        RECT 26.855 23.615 27.205 23.630 ;
        RECT 29.710 23.615 30.960 23.625 ;
        RECT 26.835 23.315 30.975 23.615 ;
        RECT 26.855 23.300 27.205 23.315 ;
        RECT 29.710 23.305 30.960 23.315 ;
        RECT 36.810 23.210 37.140 23.960 ;
        RECT 37.465 23.090 37.765 37.310 ;
        RECT 38.140 37.155 38.440 37.795 ;
        RECT 38.765 37.660 39.065 38.075 ;
        RECT 39.420 37.660 39.720 41.675 ;
        RECT 40.665 41.670 40.995 42.020 ;
        RECT 41.305 41.830 41.635 42.590 ;
        RECT 42.140 42.315 42.470 43.065 ;
        RECT 38.750 37.310 39.720 37.660 ;
        RECT 38.125 36.805 38.455 37.155 ;
        RECT 38.140 35.125 38.440 36.805 ;
        RECT 38.125 34.775 38.455 35.125 ;
        RECT 38.140 30.835 38.440 34.775 ;
        RECT 38.750 34.135 39.080 34.485 ;
        RECT 38.125 30.485 38.455 30.835 ;
        RECT 38.765 30.125 39.065 34.135 ;
        RECT 38.120 29.775 38.450 30.125 ;
        RECT 38.750 29.775 39.080 30.125 ;
        RECT 28.000 22.970 28.350 22.985 ;
        RECT 29.710 22.970 30.960 22.980 ;
        RECT 27.975 22.670 30.975 22.970 ;
        RECT 37.450 22.740 37.780 23.090 ;
        RECT 28.000 22.655 28.350 22.670 ;
        RECT 29.710 22.660 30.960 22.670 ;
        RECT 38.135 22.590 38.435 29.775 ;
        RECT 38.765 26.950 39.065 29.775 ;
        RECT 38.750 26.600 39.080 26.950 ;
        RECT 39.420 23.955 39.720 37.310 ;
        RECT 40.035 34.135 40.365 34.485 ;
        RECT 40.050 27.365 40.350 34.135 ;
        RECT 40.050 26.950 40.365 27.365 ;
        RECT 40.050 26.600 40.380 26.950 ;
        RECT 40.050 24.790 40.350 26.600 ;
        RECT 40.680 26.365 40.980 41.670 ;
        RECT 41.310 40.385 41.640 41.135 ;
        RECT 42.140 41.015 42.470 41.765 ;
        RECT 41.305 37.630 41.635 38.380 ;
        RECT 42.145 38.280 42.475 39.030 ;
        RECT 42.800 37.660 43.100 52.960 ;
        RECT 43.470 52.730 43.785 53.145 ;
        RECT 43.470 52.380 43.800 52.730 ;
        RECT 44.715 52.380 45.045 52.730 ;
        RECT 43.470 45.195 43.770 52.380 ;
        RECT 44.730 49.560 45.030 52.380 ;
        RECT 44.085 49.205 44.415 49.555 ;
        RECT 44.715 49.210 45.045 49.560 ;
        RECT 45.385 49.555 45.685 56.740 ;
        RECT 46.000 56.235 46.330 56.585 ;
        RECT 44.100 45.195 44.400 49.205 ;
        RECT 44.730 45.195 45.030 49.210 ;
        RECT 45.370 49.205 45.700 49.555 ;
        RECT 43.455 44.845 43.785 45.195 ;
        RECT 44.085 44.845 44.415 45.195 ;
        RECT 44.715 44.845 45.045 45.195 ;
        RECT 44.100 42.020 44.400 44.845 ;
        RECT 44.085 41.670 44.415 42.020 ;
        RECT 44.740 41.675 45.070 42.025 ;
        RECT 46.015 42.020 46.315 56.235 ;
        RECT 46.645 55.455 46.975 56.205 ;
        RECT 47.465 56.085 47.795 56.835 ;
        RECT 46.640 52.700 46.970 53.450 ;
        RECT 47.470 53.350 47.800 54.100 ;
        RECT 48.110 52.960 48.440 53.310 ;
        RECT 48.795 53.145 49.095 59.915 ;
        RECT 49.425 57.090 49.725 59.915 ;
        RECT 50.710 57.505 51.010 64.275 ;
        RECT 51.970 62.990 52.300 63.740 ;
        RECT 52.800 63.620 53.130 64.370 ;
        RECT 54.745 64.275 55.075 64.625 ;
        RECT 55.375 64.280 55.705 64.630 ;
        RECT 51.965 60.235 52.295 60.985 ;
        RECT 52.805 60.885 53.135 61.635 ;
        RECT 54.760 60.265 55.060 64.275 ;
        RECT 55.390 60.265 55.690 64.280 ;
        RECT 56.030 64.275 56.360 64.625 ;
        RECT 57.300 64.435 57.630 65.195 ;
        RECT 58.125 64.920 58.455 65.670 ;
        RECT 60.715 64.630 61.015 67.450 ;
        RECT 62.625 66.485 62.955 67.235 ;
        RECT 63.460 66.935 63.790 68.195 ;
        RECT 65.415 67.800 65.715 73.385 ;
        RECT 70.740 69.835 71.040 70.230 ;
        RECT 68.790 69.145 69.120 69.600 ;
        RECT 70.730 69.455 71.050 69.835 ;
        RECT 67.110 68.845 69.120 69.145 ;
        RECT 64.625 67.450 64.955 67.800 ;
        RECT 65.400 67.450 65.730 67.800 ;
        RECT 66.035 67.450 66.365 67.800 ;
        RECT 67.110 67.575 67.410 68.845 ;
        RECT 68.790 68.795 69.120 68.845 ;
        RECT 69.420 68.485 69.740 68.865 ;
        RECT 69.420 68.390 69.730 68.485 ;
        RECT 64.640 66.300 64.940 67.450 ;
        RECT 64.630 65.920 64.950 66.300 ;
        RECT 51.965 58.950 52.295 59.700 ;
        RECT 52.800 59.350 53.130 60.105 ;
        RECT 54.115 59.915 54.445 60.265 ;
        RECT 54.745 59.915 55.075 60.265 ;
        RECT 55.375 59.915 55.705 60.265 ;
        RECT 50.710 57.090 51.025 57.505 ;
        RECT 49.410 56.740 49.740 57.090 ;
        RECT 50.710 56.740 51.040 57.090 ;
        RECT 51.965 56.900 52.295 57.660 ;
        RECT 52.800 57.385 53.130 58.135 ;
        RECT 46.640 51.415 46.970 52.165 ;
        RECT 47.465 51.815 47.795 52.570 ;
        RECT 46.640 49.365 46.970 50.125 ;
        RECT 47.465 49.850 47.795 50.600 ;
        RECT 46.645 47.920 46.975 48.670 ;
        RECT 47.465 48.550 47.795 49.300 ;
        RECT 46.640 45.165 46.970 45.915 ;
        RECT 47.470 45.815 47.800 46.565 ;
        RECT 46.640 43.880 46.970 44.630 ;
        RECT 47.465 44.280 47.795 45.035 ;
        RECT 41.305 36.345 41.635 37.095 ;
        RECT 42.140 36.745 42.470 37.500 ;
        RECT 42.785 37.310 43.115 37.660 ;
        RECT 41.305 34.295 41.635 35.055 ;
        RECT 42.140 34.780 42.470 35.530 ;
        RECT 41.310 32.850 41.640 33.600 ;
        RECT 42.140 33.480 42.470 34.230 ;
        RECT 41.305 30.095 41.635 30.845 ;
        RECT 42.145 30.745 42.475 31.495 ;
        RECT 41.305 28.810 41.635 29.560 ;
        RECT 42.140 29.210 42.470 29.965 ;
        RECT 41.305 26.760 41.635 27.520 ;
        RECT 42.140 27.245 42.470 27.995 ;
        RECT 40.665 26.015 40.995 26.365 ;
        RECT 41.310 25.315 41.640 26.065 ;
        RECT 42.140 25.945 42.470 26.695 ;
        RECT 40.050 24.490 40.990 24.790 ;
        RECT 39.420 23.655 40.355 23.955 ;
        RECT 26.480 22.325 26.830 22.340 ;
        RECT 29.710 22.325 30.960 22.335 ;
        RECT 26.460 22.025 30.975 22.325 ;
        RECT 26.480 22.010 26.830 22.025 ;
        RECT 29.710 22.015 30.960 22.025 ;
        RECT 28.380 21.680 28.730 21.695 ;
        RECT 29.710 21.680 30.960 21.690 ;
        RECT 28.340 21.380 30.975 21.680 ;
        RECT 36.805 21.675 37.135 22.430 ;
        RECT 38.120 22.240 38.450 22.590 ;
        RECT 39.380 22.240 39.710 22.590 ;
        RECT 28.380 21.365 28.730 21.380 ;
        RECT 29.710 21.370 30.960 21.380 ;
        RECT 27.995 20.350 28.345 20.365 ;
        RECT 27.995 20.345 28.760 20.350 ;
        RECT 29.710 20.345 30.960 20.355 ;
        RECT 27.975 20.045 30.975 20.345 ;
        RECT 27.995 20.035 28.345 20.045 ;
        RECT 29.710 20.035 30.960 20.045 ;
        RECT 27.620 19.700 27.970 19.715 ;
        RECT 36.805 19.710 37.135 20.460 ;
        RECT 29.710 19.700 30.960 19.710 ;
        RECT 27.620 19.400 30.975 19.700 ;
        RECT 27.620 19.385 27.970 19.400 ;
        RECT 29.710 19.390 30.960 19.400 ;
        RECT 28.380 19.055 28.730 19.070 ;
        RECT 29.710 19.055 30.960 19.065 ;
        RECT 28.355 18.755 30.975 19.055 ;
        RECT 28.380 18.740 28.730 18.755 ;
        RECT 29.710 18.745 30.960 18.755 ;
        RECT 27.240 18.410 27.590 18.425 ;
        RECT 29.710 18.410 30.960 18.420 ;
        RECT 36.805 18.410 37.135 19.160 ;
        RECT 27.215 18.110 30.975 18.410 ;
        RECT 27.240 18.095 27.590 18.110 ;
        RECT 29.710 18.100 30.960 18.110 ;
        RECT 27.615 16.080 27.965 16.095 ;
        RECT 29.710 16.080 30.960 16.090 ;
        RECT 27.615 15.780 30.975 16.080 ;
        RECT 27.615 15.765 27.965 15.780 ;
        RECT 29.710 15.770 30.960 15.780 ;
        RECT 36.810 15.675 37.140 16.425 ;
        RECT 28.380 15.435 28.730 15.450 ;
        RECT 29.710 15.435 30.960 15.445 ;
        RECT 28.370 15.135 30.975 15.435 ;
        RECT 28.380 15.120 28.730 15.135 ;
        RECT 29.710 15.125 30.960 15.135 ;
        RECT 38.135 15.055 38.435 22.240 ;
        RECT 39.395 19.420 39.695 22.240 ;
        RECT 38.750 19.065 39.080 19.415 ;
        RECT 39.380 19.070 39.710 19.420 ;
        RECT 38.765 15.055 39.065 19.065 ;
        RECT 39.395 15.055 39.695 19.070 ;
        RECT 27.240 14.790 27.590 14.805 ;
        RECT 29.710 14.790 30.960 14.800 ;
        RECT 27.195 14.490 30.975 14.790 ;
        RECT 27.240 14.475 27.590 14.490 ;
        RECT 29.710 14.480 30.960 14.490 ;
        RECT 28.000 14.145 28.350 14.160 ;
        RECT 29.710 14.145 30.960 14.155 ;
        RECT 27.985 13.845 30.975 14.145 ;
        RECT 36.805 14.140 37.135 14.895 ;
        RECT 38.120 14.705 38.450 15.055 ;
        RECT 38.750 14.705 39.080 15.055 ;
        RECT 39.380 14.705 39.710 15.055 ;
        RECT 28.000 13.830 28.350 13.845 ;
        RECT 29.710 13.835 30.960 13.845 ;
        RECT 28.375 12.810 28.725 12.825 ;
        RECT 29.710 12.810 30.960 12.820 ;
        RECT 28.325 12.510 30.975 12.810 ;
        RECT 28.375 12.495 28.725 12.510 ;
        RECT 29.710 12.500 30.960 12.510 ;
        RECT 24.960 12.165 25.310 12.180 ;
        RECT 36.805 12.175 37.135 12.925 ;
        RECT 29.710 12.165 30.960 12.175 ;
        RECT 24.960 11.865 30.975 12.165 ;
        RECT 38.765 11.880 39.065 14.705 ;
        RECT 24.960 11.850 25.310 11.865 ;
        RECT 29.710 11.855 30.960 11.865 ;
        RECT 28.000 11.520 28.350 11.530 ;
        RECT 29.710 11.520 30.960 11.530 ;
        RECT 27.990 11.220 30.975 11.520 ;
        RECT 28.000 11.215 28.765 11.220 ;
        RECT 28.000 11.200 28.350 11.215 ;
        RECT 29.710 11.210 30.960 11.220 ;
        RECT 25.340 10.875 25.690 10.890 ;
        RECT 29.710 10.875 30.960 10.885 ;
        RECT 36.805 10.875 37.135 11.625 ;
        RECT 38.750 11.530 39.080 11.880 ;
        RECT 39.390 11.535 39.720 11.885 ;
        RECT 40.055 11.880 40.355 23.655 ;
        RECT 40.690 19.415 40.990 24.490 ;
        RECT 41.305 22.560 41.635 23.310 ;
        RECT 42.145 23.210 42.475 23.960 ;
        RECT 42.800 23.090 43.100 37.310 ;
        RECT 43.475 37.155 43.775 37.795 ;
        RECT 44.100 37.660 44.400 38.075 ;
        RECT 44.755 37.660 45.055 41.675 ;
        RECT 46.000 41.670 46.330 42.020 ;
        RECT 46.640 41.830 46.970 42.590 ;
        RECT 47.465 42.315 47.795 43.065 ;
        RECT 44.085 37.310 45.055 37.660 ;
        RECT 43.460 36.805 43.790 37.155 ;
        RECT 43.475 35.125 43.775 36.805 ;
        RECT 43.460 34.775 43.790 35.125 ;
        RECT 43.475 30.835 43.775 34.775 ;
        RECT 44.085 34.135 44.415 34.485 ;
        RECT 43.460 30.485 43.790 30.835 ;
        RECT 44.100 30.125 44.400 34.135 ;
        RECT 43.455 29.775 43.785 30.125 ;
        RECT 44.085 29.775 44.415 30.125 ;
        RECT 42.785 22.740 43.115 23.090 ;
        RECT 43.470 22.590 43.770 29.775 ;
        RECT 44.100 26.950 44.400 29.775 ;
        RECT 44.085 26.600 44.415 26.950 ;
        RECT 44.755 23.955 45.055 37.310 ;
        RECT 45.370 34.135 45.700 34.485 ;
        RECT 45.385 27.365 45.685 34.135 ;
        RECT 45.385 26.950 45.700 27.365 ;
        RECT 45.385 26.600 45.715 26.950 ;
        RECT 45.385 24.790 45.685 26.600 ;
        RECT 46.015 26.365 46.315 41.670 ;
        RECT 46.645 40.385 46.975 41.135 ;
        RECT 47.465 41.015 47.795 41.765 ;
        RECT 46.640 37.630 46.970 38.380 ;
        RECT 47.470 38.280 47.800 39.030 ;
        RECT 48.125 37.660 48.425 52.960 ;
        RECT 48.795 52.730 49.110 53.145 ;
        RECT 48.795 52.380 49.125 52.730 ;
        RECT 50.040 52.380 50.370 52.730 ;
        RECT 48.795 45.195 49.095 52.380 ;
        RECT 50.055 49.560 50.355 52.380 ;
        RECT 49.410 49.205 49.740 49.555 ;
        RECT 50.040 49.210 50.370 49.560 ;
        RECT 50.710 49.555 51.010 56.740 ;
        RECT 51.325 56.235 51.655 56.585 ;
        RECT 49.425 45.195 49.725 49.205 ;
        RECT 50.055 45.195 50.355 49.210 ;
        RECT 50.695 49.205 51.025 49.555 ;
        RECT 48.780 44.845 49.110 45.195 ;
        RECT 49.410 44.845 49.740 45.195 ;
        RECT 50.040 44.845 50.370 45.195 ;
        RECT 49.425 42.020 49.725 44.845 ;
        RECT 49.410 41.670 49.740 42.020 ;
        RECT 50.065 41.675 50.395 42.025 ;
        RECT 51.340 42.020 51.640 56.235 ;
        RECT 51.970 55.455 52.300 56.205 ;
        RECT 52.800 56.085 53.130 56.835 ;
        RECT 51.965 52.700 52.295 53.450 ;
        RECT 52.805 53.350 53.135 54.100 ;
        RECT 53.445 52.960 53.775 53.310 ;
        RECT 54.130 53.145 54.430 59.915 ;
        RECT 54.760 57.090 55.060 59.915 ;
        RECT 56.045 57.505 56.345 64.275 ;
        RECT 57.305 62.990 57.635 63.740 ;
        RECT 58.125 63.620 58.455 64.370 ;
        RECT 60.070 64.275 60.400 64.625 ;
        RECT 60.700 64.280 61.030 64.630 ;
        RECT 57.300 60.235 57.630 60.985 ;
        RECT 58.130 60.885 58.460 61.635 ;
        RECT 60.085 60.265 60.385 64.275 ;
        RECT 60.715 60.265 61.015 64.280 ;
        RECT 61.355 64.275 61.685 64.625 ;
        RECT 62.625 64.435 62.955 65.195 ;
        RECT 63.460 64.920 63.790 65.670 ;
        RECT 66.050 64.630 66.350 67.450 ;
        RECT 67.100 67.195 67.420 67.575 ;
        RECT 67.960 67.535 68.290 68.270 ;
        RECT 68.785 68.090 69.730 68.390 ;
        RECT 67.960 66.485 68.290 67.235 ;
        RECT 68.785 66.935 69.115 68.090 ;
        RECT 70.740 67.800 71.040 69.455 ;
        RECT 69.950 67.450 70.280 67.800 ;
        RECT 70.725 67.450 71.055 67.800 ;
        RECT 71.360 67.450 71.690 67.800 ;
        RECT 73.285 67.535 73.615 68.270 ;
        RECT 76.075 67.800 76.375 70.185 ;
        RECT 81.400 69.835 81.700 70.230 ;
        RECT 79.450 68.795 79.780 69.600 ;
        RECT 81.390 69.455 81.710 69.835 ;
        RECT 85.450 69.820 85.750 79.750 ;
        RECT 86.080 79.710 86.380 80.125 ;
        RECT 86.065 79.360 86.395 79.710 ;
        RECT 84.785 69.520 85.750 69.820 ;
        RECT 79.450 68.485 79.770 68.795 ;
        RECT 75.285 67.450 75.615 67.800 ;
        RECT 76.060 67.450 76.390 67.800 ;
        RECT 76.695 67.450 77.025 67.800 ;
        RECT 78.620 67.535 78.950 68.270 ;
        RECT 79.460 67.670 79.760 67.970 ;
        RECT 81.400 67.800 81.700 69.455 ;
        RECT 84.785 68.795 85.115 69.520 ;
        RECT 86.080 68.495 86.380 79.360 ;
        RECT 86.725 73.385 87.045 73.765 ;
        RECT 69.965 66.300 70.265 67.450 ;
        RECT 69.955 65.920 70.275 66.300 ;
        RECT 57.300 58.950 57.630 59.700 ;
        RECT 58.125 59.350 58.455 60.105 ;
        RECT 59.440 59.915 59.770 60.265 ;
        RECT 60.070 59.915 60.400 60.265 ;
        RECT 60.700 59.915 61.030 60.265 ;
        RECT 56.045 57.090 56.360 57.505 ;
        RECT 54.745 56.740 55.075 57.090 ;
        RECT 56.045 56.740 56.375 57.090 ;
        RECT 57.300 56.900 57.630 57.660 ;
        RECT 58.125 57.385 58.455 58.135 ;
        RECT 51.965 51.415 52.295 52.165 ;
        RECT 52.800 51.815 53.130 52.570 ;
        RECT 51.965 49.365 52.295 50.125 ;
        RECT 52.800 49.850 53.130 50.600 ;
        RECT 51.970 47.920 52.300 48.670 ;
        RECT 52.800 48.550 53.130 49.300 ;
        RECT 51.965 45.165 52.295 45.915 ;
        RECT 52.805 45.815 53.135 46.565 ;
        RECT 51.965 43.880 52.295 44.630 ;
        RECT 52.800 44.280 53.130 45.035 ;
        RECT 46.640 36.345 46.970 37.095 ;
        RECT 47.465 36.745 47.795 37.500 ;
        RECT 48.110 37.310 48.440 37.660 ;
        RECT 46.640 34.295 46.970 35.055 ;
        RECT 47.465 34.780 47.795 35.530 ;
        RECT 46.645 32.850 46.975 33.600 ;
        RECT 47.465 33.480 47.795 34.230 ;
        RECT 46.640 30.095 46.970 30.845 ;
        RECT 47.470 30.745 47.800 31.495 ;
        RECT 46.640 28.810 46.970 29.560 ;
        RECT 47.465 29.210 47.795 29.965 ;
        RECT 46.640 26.760 46.970 27.520 ;
        RECT 47.465 27.245 47.795 27.995 ;
        RECT 46.000 26.015 46.330 26.365 ;
        RECT 46.645 25.315 46.975 26.065 ;
        RECT 47.465 25.945 47.795 26.695 ;
        RECT 45.385 24.490 46.325 24.790 ;
        RECT 44.755 23.655 45.690 23.955 ;
        RECT 41.305 21.275 41.635 22.025 ;
        RECT 42.140 21.675 42.470 22.430 ;
        RECT 43.455 22.240 43.785 22.590 ;
        RECT 44.715 22.240 45.045 22.590 ;
        RECT 40.675 19.065 41.005 19.415 ;
        RECT 41.305 19.225 41.635 19.985 ;
        RECT 42.140 19.710 42.470 20.460 ;
        RECT 41.310 17.780 41.640 18.530 ;
        RECT 42.140 18.410 42.470 19.160 ;
        RECT 41.305 15.025 41.635 15.775 ;
        RECT 42.145 15.675 42.475 16.425 ;
        RECT 43.470 15.055 43.770 22.240 ;
        RECT 44.730 19.420 45.030 22.240 ;
        RECT 44.085 19.065 44.415 19.415 ;
        RECT 44.715 19.070 45.045 19.420 ;
        RECT 44.100 15.055 44.400 19.065 ;
        RECT 44.730 15.055 45.030 19.070 ;
        RECT 41.305 13.740 41.635 14.490 ;
        RECT 42.140 14.140 42.470 14.895 ;
        RECT 43.455 14.705 43.785 15.055 ;
        RECT 44.085 14.705 44.415 15.055 ;
        RECT 44.715 14.705 45.045 15.055 ;
        RECT 25.340 10.575 30.975 10.875 ;
        RECT 25.340 10.560 25.690 10.575 ;
        RECT 29.710 10.565 30.960 10.575 ;
        RECT 39.405 9.590 39.705 11.535 ;
        RECT 40.040 11.530 40.370 11.880 ;
        RECT 41.305 11.690 41.635 12.450 ;
        RECT 42.140 12.175 42.470 12.925 ;
        RECT 44.100 11.880 44.400 14.705 ;
        RECT 41.310 10.245 41.640 10.995 ;
        RECT 42.140 10.875 42.470 11.625 ;
        RECT 44.085 11.530 44.415 11.880 ;
        RECT 44.725 11.535 45.055 11.885 ;
        RECT 45.390 11.880 45.690 23.655 ;
        RECT 46.025 19.415 46.325 24.490 ;
        RECT 46.640 22.560 46.970 23.310 ;
        RECT 47.470 23.210 47.800 23.960 ;
        RECT 48.125 23.090 48.425 37.310 ;
        RECT 48.800 37.155 49.100 37.795 ;
        RECT 49.425 37.660 49.725 38.075 ;
        RECT 50.080 37.660 50.380 41.675 ;
        RECT 51.325 41.670 51.655 42.020 ;
        RECT 51.965 41.830 52.295 42.590 ;
        RECT 52.800 42.315 53.130 43.065 ;
        RECT 49.410 37.310 50.380 37.660 ;
        RECT 48.785 36.805 49.115 37.155 ;
        RECT 48.800 35.125 49.100 36.805 ;
        RECT 48.785 34.775 49.115 35.125 ;
        RECT 48.800 30.835 49.100 34.775 ;
        RECT 49.410 34.135 49.740 34.485 ;
        RECT 48.785 30.485 49.115 30.835 ;
        RECT 49.425 30.125 49.725 34.135 ;
        RECT 48.780 29.775 49.110 30.125 ;
        RECT 49.410 29.775 49.740 30.125 ;
        RECT 48.110 22.740 48.440 23.090 ;
        RECT 48.795 22.590 49.095 29.775 ;
        RECT 49.425 26.950 49.725 29.775 ;
        RECT 49.410 26.600 49.740 26.950 ;
        RECT 50.080 23.955 50.380 37.310 ;
        RECT 50.695 34.135 51.025 34.485 ;
        RECT 50.710 27.365 51.010 34.135 ;
        RECT 50.710 26.950 51.025 27.365 ;
        RECT 50.710 26.600 51.040 26.950 ;
        RECT 50.710 24.790 51.010 26.600 ;
        RECT 51.340 26.365 51.640 41.670 ;
        RECT 51.970 40.385 52.300 41.135 ;
        RECT 52.800 41.015 53.130 41.765 ;
        RECT 51.965 37.630 52.295 38.380 ;
        RECT 52.805 38.280 53.135 39.030 ;
        RECT 53.460 37.660 53.760 52.960 ;
        RECT 54.130 52.730 54.445 53.145 ;
        RECT 54.130 52.380 54.460 52.730 ;
        RECT 55.375 52.380 55.705 52.730 ;
        RECT 54.130 45.195 54.430 52.380 ;
        RECT 55.390 49.560 55.690 52.380 ;
        RECT 54.745 49.205 55.075 49.555 ;
        RECT 55.375 49.210 55.705 49.560 ;
        RECT 56.045 49.555 56.345 56.740 ;
        RECT 56.660 56.235 56.990 56.585 ;
        RECT 54.760 45.195 55.060 49.205 ;
        RECT 55.390 45.195 55.690 49.210 ;
        RECT 56.030 49.205 56.360 49.555 ;
        RECT 54.115 44.845 54.445 45.195 ;
        RECT 54.745 44.845 55.075 45.195 ;
        RECT 55.375 44.845 55.705 45.195 ;
        RECT 54.760 42.020 55.060 44.845 ;
        RECT 54.745 41.670 55.075 42.020 ;
        RECT 55.400 41.675 55.730 42.025 ;
        RECT 56.675 42.020 56.975 56.235 ;
        RECT 57.305 55.455 57.635 56.205 ;
        RECT 58.125 56.085 58.455 56.835 ;
        RECT 57.300 52.700 57.630 53.450 ;
        RECT 58.130 53.350 58.460 54.100 ;
        RECT 58.770 52.960 59.100 53.310 ;
        RECT 59.455 53.145 59.755 59.915 ;
        RECT 60.085 57.090 60.385 59.915 ;
        RECT 61.370 57.505 61.670 64.275 ;
        RECT 62.630 62.990 62.960 63.740 ;
        RECT 63.460 63.620 63.790 64.370 ;
        RECT 65.405 64.275 65.735 64.625 ;
        RECT 66.035 64.280 66.365 64.630 ;
        RECT 62.625 60.235 62.955 60.985 ;
        RECT 63.465 60.885 63.795 61.635 ;
        RECT 65.420 60.265 65.720 64.275 ;
        RECT 66.050 60.265 66.350 64.280 ;
        RECT 66.690 64.275 67.020 64.625 ;
        RECT 67.960 64.435 68.290 65.195 ;
        RECT 68.785 64.920 69.115 65.670 ;
        RECT 71.375 64.630 71.675 67.450 ;
        RECT 73.285 66.485 73.615 67.235 ;
        RECT 75.300 66.300 75.600 67.450 ;
        RECT 75.290 65.920 75.610 66.300 ;
        RECT 62.625 58.950 62.955 59.700 ;
        RECT 63.460 59.350 63.790 60.105 ;
        RECT 64.775 59.915 65.105 60.265 ;
        RECT 65.405 59.915 65.735 60.265 ;
        RECT 66.035 59.915 66.365 60.265 ;
        RECT 61.370 57.090 61.685 57.505 ;
        RECT 60.070 56.740 60.400 57.090 ;
        RECT 61.370 56.740 61.700 57.090 ;
        RECT 62.625 56.900 62.955 57.660 ;
        RECT 63.460 57.385 63.790 58.135 ;
        RECT 57.300 51.415 57.630 52.165 ;
        RECT 58.125 51.815 58.455 52.570 ;
        RECT 57.300 49.365 57.630 50.125 ;
        RECT 58.125 49.850 58.455 50.600 ;
        RECT 57.305 47.920 57.635 48.670 ;
        RECT 58.125 48.550 58.455 49.300 ;
        RECT 57.300 45.165 57.630 45.915 ;
        RECT 58.130 45.815 58.460 46.565 ;
        RECT 57.300 43.880 57.630 44.630 ;
        RECT 58.125 44.280 58.455 45.035 ;
        RECT 51.965 36.345 52.295 37.095 ;
        RECT 52.800 36.745 53.130 37.500 ;
        RECT 53.445 37.310 53.775 37.660 ;
        RECT 51.965 34.295 52.295 35.055 ;
        RECT 52.800 34.780 53.130 35.530 ;
        RECT 51.970 32.850 52.300 33.600 ;
        RECT 52.800 33.480 53.130 34.230 ;
        RECT 51.965 30.095 52.295 30.845 ;
        RECT 52.805 30.745 53.135 31.495 ;
        RECT 51.965 28.810 52.295 29.560 ;
        RECT 52.800 29.210 53.130 29.965 ;
        RECT 51.965 26.760 52.295 27.520 ;
        RECT 52.800 27.245 53.130 27.995 ;
        RECT 51.325 26.015 51.655 26.365 ;
        RECT 51.970 25.315 52.300 26.065 ;
        RECT 52.800 25.945 53.130 26.695 ;
        RECT 50.710 24.490 51.650 24.790 ;
        RECT 50.080 23.655 51.015 23.955 ;
        RECT 46.640 21.275 46.970 22.025 ;
        RECT 47.465 21.675 47.795 22.430 ;
        RECT 48.780 22.240 49.110 22.590 ;
        RECT 50.040 22.240 50.370 22.590 ;
        RECT 46.010 19.065 46.340 19.415 ;
        RECT 46.640 19.225 46.970 19.985 ;
        RECT 47.465 19.710 47.795 20.460 ;
        RECT 46.645 17.780 46.975 18.530 ;
        RECT 47.465 18.410 47.795 19.160 ;
        RECT 46.640 15.025 46.970 15.775 ;
        RECT 47.470 15.675 47.800 16.425 ;
        RECT 48.795 15.055 49.095 22.240 ;
        RECT 50.055 19.420 50.355 22.240 ;
        RECT 49.410 19.065 49.740 19.415 ;
        RECT 50.040 19.070 50.370 19.420 ;
        RECT 49.425 15.055 49.725 19.065 ;
        RECT 50.055 15.055 50.355 19.070 ;
        RECT 46.640 13.740 46.970 14.490 ;
        RECT 47.465 14.140 47.795 14.895 ;
        RECT 48.780 14.705 49.110 15.055 ;
        RECT 49.410 14.705 49.740 15.055 ;
        RECT 50.040 14.705 50.370 15.055 ;
        RECT 44.740 9.750 45.040 11.535 ;
        RECT 45.375 11.530 45.705 11.880 ;
        RECT 46.640 11.620 46.970 12.450 ;
        RECT 47.465 12.175 47.795 12.925 ;
        RECT 49.425 11.880 49.725 14.705 ;
        RECT 46.020 11.310 46.970 11.620 ;
        RECT 46.020 10.610 46.330 11.310 ;
        RECT 46.010 10.240 46.340 10.610 ;
        RECT 46.645 10.245 46.975 10.995 ;
        RECT 47.465 10.875 47.795 11.625 ;
        RECT 49.410 11.530 49.740 11.880 ;
        RECT 50.050 11.535 50.380 11.885 ;
        RECT 50.715 11.880 51.015 23.655 ;
        RECT 51.350 19.415 51.650 24.490 ;
        RECT 51.965 22.560 52.295 23.310 ;
        RECT 52.805 23.210 53.135 23.960 ;
        RECT 53.460 23.090 53.760 37.310 ;
        RECT 54.135 37.155 54.435 37.795 ;
        RECT 54.760 37.660 55.060 38.075 ;
        RECT 55.415 37.660 55.715 41.675 ;
        RECT 56.660 41.670 56.990 42.020 ;
        RECT 57.300 41.830 57.630 42.590 ;
        RECT 58.125 42.315 58.455 43.065 ;
        RECT 54.745 37.310 55.715 37.660 ;
        RECT 54.120 36.805 54.450 37.155 ;
        RECT 54.135 35.125 54.435 36.805 ;
        RECT 54.120 34.775 54.450 35.125 ;
        RECT 54.135 30.835 54.435 34.775 ;
        RECT 54.745 34.135 55.075 34.485 ;
        RECT 54.120 30.485 54.450 30.835 ;
        RECT 54.760 30.125 55.060 34.135 ;
        RECT 54.115 29.775 54.445 30.125 ;
        RECT 54.745 29.775 55.075 30.125 ;
        RECT 53.445 22.740 53.775 23.090 ;
        RECT 54.130 22.590 54.430 29.775 ;
        RECT 54.760 26.950 55.060 29.775 ;
        RECT 54.745 26.600 55.075 26.950 ;
        RECT 55.415 23.955 55.715 37.310 ;
        RECT 56.030 34.135 56.360 34.485 ;
        RECT 56.045 27.365 56.345 34.135 ;
        RECT 56.045 26.950 56.360 27.365 ;
        RECT 56.045 26.600 56.375 26.950 ;
        RECT 56.045 24.790 56.345 26.600 ;
        RECT 56.675 26.365 56.975 41.670 ;
        RECT 57.305 40.385 57.635 41.135 ;
        RECT 58.125 41.015 58.455 41.765 ;
        RECT 57.300 37.630 57.630 38.380 ;
        RECT 58.130 38.280 58.460 39.030 ;
        RECT 58.785 37.660 59.085 52.960 ;
        RECT 59.455 52.730 59.770 53.145 ;
        RECT 59.455 52.380 59.785 52.730 ;
        RECT 60.700 52.380 61.030 52.730 ;
        RECT 59.455 45.195 59.755 52.380 ;
        RECT 60.715 49.560 61.015 52.380 ;
        RECT 60.070 49.205 60.400 49.555 ;
        RECT 60.700 49.210 61.030 49.560 ;
        RECT 61.370 49.555 61.670 56.740 ;
        RECT 61.985 56.235 62.315 56.585 ;
        RECT 60.085 45.195 60.385 49.205 ;
        RECT 60.715 45.195 61.015 49.210 ;
        RECT 61.355 49.205 61.685 49.555 ;
        RECT 59.440 44.845 59.770 45.195 ;
        RECT 60.070 44.845 60.400 45.195 ;
        RECT 60.700 44.845 61.030 45.195 ;
        RECT 60.085 42.020 60.385 44.845 ;
        RECT 60.070 41.670 60.400 42.020 ;
        RECT 60.725 41.675 61.055 42.025 ;
        RECT 62.000 42.020 62.300 56.235 ;
        RECT 62.630 55.455 62.960 56.205 ;
        RECT 63.460 56.085 63.790 56.835 ;
        RECT 62.625 52.700 62.955 53.450 ;
        RECT 63.465 53.350 63.795 54.100 ;
        RECT 64.105 52.960 64.435 53.310 ;
        RECT 64.790 53.145 65.090 59.915 ;
        RECT 65.420 57.090 65.720 59.915 ;
        RECT 66.705 57.505 67.005 64.275 ;
        RECT 67.965 62.990 68.295 63.740 ;
        RECT 68.785 63.620 69.115 64.370 ;
        RECT 70.730 64.275 71.060 64.625 ;
        RECT 71.360 64.280 71.690 64.630 ;
        RECT 67.960 60.235 68.290 60.985 ;
        RECT 68.790 60.885 69.120 61.635 ;
        RECT 70.745 60.265 71.045 64.275 ;
        RECT 71.375 60.265 71.675 64.280 ;
        RECT 72.015 64.275 72.345 64.625 ;
        RECT 73.285 64.435 73.615 65.195 ;
        RECT 74.120 64.920 74.450 65.670 ;
        RECT 76.710 64.630 77.010 67.450 ;
        RECT 77.600 66.300 77.900 66.695 ;
        RECT 78.620 66.485 78.950 67.235 ;
        RECT 79.445 66.935 79.775 67.670 ;
        RECT 80.610 67.450 80.940 67.800 ;
        RECT 81.385 67.450 81.715 67.800 ;
        RECT 82.020 67.450 82.350 67.800 ;
        RECT 83.945 67.535 84.275 68.270 ;
        RECT 84.780 68.195 86.380 68.495 ;
        RECT 80.625 66.300 80.925 67.450 ;
        RECT 77.590 65.920 77.910 66.300 ;
        RECT 80.615 65.920 80.935 66.300 ;
        RECT 67.960 58.950 68.290 59.700 ;
        RECT 68.785 59.350 69.115 60.105 ;
        RECT 70.100 59.915 70.430 60.265 ;
        RECT 70.730 59.915 71.060 60.265 ;
        RECT 71.360 59.915 71.690 60.265 ;
        RECT 66.705 57.090 67.020 57.505 ;
        RECT 65.405 56.740 65.735 57.090 ;
        RECT 66.705 56.740 67.035 57.090 ;
        RECT 67.960 56.900 68.290 57.660 ;
        RECT 68.785 57.385 69.115 58.135 ;
        RECT 62.625 51.415 62.955 52.165 ;
        RECT 63.460 51.815 63.790 52.570 ;
        RECT 62.625 49.365 62.955 50.125 ;
        RECT 63.460 49.850 63.790 50.600 ;
        RECT 62.630 47.920 62.960 48.670 ;
        RECT 63.460 48.550 63.790 49.300 ;
        RECT 62.625 45.165 62.955 45.915 ;
        RECT 63.465 45.815 63.795 46.565 ;
        RECT 62.625 43.880 62.955 44.630 ;
        RECT 63.460 44.280 63.790 45.035 ;
        RECT 57.300 36.345 57.630 37.095 ;
        RECT 58.125 36.745 58.455 37.500 ;
        RECT 58.770 37.310 59.100 37.660 ;
        RECT 57.300 34.295 57.630 35.055 ;
        RECT 58.125 34.780 58.455 35.530 ;
        RECT 57.305 32.850 57.635 33.600 ;
        RECT 58.125 33.480 58.455 34.230 ;
        RECT 57.300 30.095 57.630 30.845 ;
        RECT 58.130 30.745 58.460 31.495 ;
        RECT 57.300 28.810 57.630 29.560 ;
        RECT 58.125 29.210 58.455 29.965 ;
        RECT 57.300 26.760 57.630 27.520 ;
        RECT 58.125 27.245 58.455 27.995 ;
        RECT 56.660 26.015 56.990 26.365 ;
        RECT 57.305 25.315 57.635 26.065 ;
        RECT 58.125 25.945 58.455 26.695 ;
        RECT 56.045 24.490 56.985 24.790 ;
        RECT 55.415 23.655 56.350 23.955 ;
        RECT 51.965 21.275 52.295 22.025 ;
        RECT 52.800 21.675 53.130 22.430 ;
        RECT 54.115 22.240 54.445 22.590 ;
        RECT 55.375 22.240 55.705 22.590 ;
        RECT 51.335 19.065 51.665 19.415 ;
        RECT 51.965 19.225 52.295 19.985 ;
        RECT 52.800 19.710 53.130 20.460 ;
        RECT 51.970 17.780 52.300 18.530 ;
        RECT 52.800 18.410 53.130 19.160 ;
        RECT 51.965 15.025 52.295 15.775 ;
        RECT 52.805 15.675 53.135 16.425 ;
        RECT 54.130 15.055 54.430 22.240 ;
        RECT 55.390 19.420 55.690 22.240 ;
        RECT 54.745 19.065 55.075 19.415 ;
        RECT 55.375 19.070 55.705 19.420 ;
        RECT 54.760 15.055 55.060 19.065 ;
        RECT 55.390 15.055 55.690 19.070 ;
        RECT 51.965 13.740 52.295 14.490 ;
        RECT 52.800 14.140 53.130 14.895 ;
        RECT 54.115 14.705 54.445 15.055 ;
        RECT 54.745 14.705 55.075 15.055 ;
        RECT 55.375 14.705 55.705 15.055 ;
        RECT 39.395 9.210 39.715 9.590 ;
        RECT 44.730 9.370 45.050 9.750 ;
        RECT 50.065 9.590 50.365 11.535 ;
        RECT 50.700 11.530 51.030 11.880 ;
        RECT 51.965 11.690 52.295 12.450 ;
        RECT 52.800 12.175 53.130 12.925 ;
        RECT 54.760 11.880 55.060 14.705 ;
        RECT 51.970 10.245 52.300 10.995 ;
        RECT 52.800 10.875 53.130 11.625 ;
        RECT 54.745 11.530 55.075 11.880 ;
        RECT 55.385 11.535 55.715 11.885 ;
        RECT 56.050 11.880 56.350 23.655 ;
        RECT 56.685 19.415 56.985 24.490 ;
        RECT 57.300 22.560 57.630 23.310 ;
        RECT 58.130 23.210 58.460 23.960 ;
        RECT 58.785 23.090 59.085 37.310 ;
        RECT 59.460 37.155 59.760 37.795 ;
        RECT 60.085 37.660 60.385 38.075 ;
        RECT 60.740 37.660 61.040 41.675 ;
        RECT 61.985 41.670 62.315 42.020 ;
        RECT 62.625 41.830 62.955 42.590 ;
        RECT 63.460 42.315 63.790 43.065 ;
        RECT 60.070 37.310 61.040 37.660 ;
        RECT 59.445 36.805 59.775 37.155 ;
        RECT 59.460 35.125 59.760 36.805 ;
        RECT 59.445 34.775 59.775 35.125 ;
        RECT 59.460 30.835 59.760 34.775 ;
        RECT 60.070 34.135 60.400 34.485 ;
        RECT 59.445 30.485 59.775 30.835 ;
        RECT 60.085 30.125 60.385 34.135 ;
        RECT 59.440 29.775 59.770 30.125 ;
        RECT 60.070 29.775 60.400 30.125 ;
        RECT 58.770 22.740 59.100 23.090 ;
        RECT 59.455 22.590 59.755 29.775 ;
        RECT 60.085 26.950 60.385 29.775 ;
        RECT 60.070 26.600 60.400 26.950 ;
        RECT 60.740 23.955 61.040 37.310 ;
        RECT 61.355 34.135 61.685 34.485 ;
        RECT 61.370 27.365 61.670 34.135 ;
        RECT 61.370 26.950 61.685 27.365 ;
        RECT 61.370 26.600 61.700 26.950 ;
        RECT 61.370 24.790 61.670 26.600 ;
        RECT 62.000 26.365 62.300 41.670 ;
        RECT 62.630 40.385 62.960 41.135 ;
        RECT 63.460 41.015 63.790 41.765 ;
        RECT 62.625 37.630 62.955 38.380 ;
        RECT 63.465 38.280 63.795 39.030 ;
        RECT 64.120 37.660 64.420 52.960 ;
        RECT 64.790 52.730 65.105 53.145 ;
        RECT 64.790 52.380 65.120 52.730 ;
        RECT 66.035 52.380 66.365 52.730 ;
        RECT 64.790 45.195 65.090 52.380 ;
        RECT 66.050 49.560 66.350 52.380 ;
        RECT 65.405 49.205 65.735 49.555 ;
        RECT 66.035 49.210 66.365 49.560 ;
        RECT 66.705 49.555 67.005 56.740 ;
        RECT 67.320 56.235 67.650 56.585 ;
        RECT 65.420 45.195 65.720 49.205 ;
        RECT 66.050 45.195 66.350 49.210 ;
        RECT 66.690 49.205 67.020 49.555 ;
        RECT 64.775 44.845 65.105 45.195 ;
        RECT 65.405 44.845 65.735 45.195 ;
        RECT 66.035 44.845 66.365 45.195 ;
        RECT 65.420 42.020 65.720 44.845 ;
        RECT 65.405 41.670 65.735 42.020 ;
        RECT 66.060 41.675 66.390 42.025 ;
        RECT 67.335 42.020 67.635 56.235 ;
        RECT 67.965 55.455 68.295 56.205 ;
        RECT 68.785 56.085 69.115 56.835 ;
        RECT 67.960 52.700 68.290 53.450 ;
        RECT 68.790 53.350 69.120 54.100 ;
        RECT 69.430 52.960 69.760 53.310 ;
        RECT 70.115 53.145 70.415 59.915 ;
        RECT 70.745 57.090 71.045 59.915 ;
        RECT 72.030 57.505 72.330 64.275 ;
        RECT 73.290 62.990 73.620 63.740 ;
        RECT 74.120 63.620 74.450 64.370 ;
        RECT 76.065 64.275 76.395 64.625 ;
        RECT 76.695 64.280 77.025 64.630 ;
        RECT 73.285 60.235 73.615 60.985 ;
        RECT 74.125 60.885 74.455 61.635 ;
        RECT 76.080 60.265 76.380 64.275 ;
        RECT 76.710 60.265 77.010 64.280 ;
        RECT 77.350 64.275 77.680 64.625 ;
        RECT 78.620 64.435 78.950 65.195 ;
        RECT 79.445 64.920 79.775 65.670 ;
        RECT 82.035 64.630 82.335 67.450 ;
        RECT 83.945 66.485 84.275 67.235 ;
        RECT 84.780 66.935 85.110 68.195 ;
        RECT 86.735 67.800 87.035 73.385 ;
        RECT 92.060 69.835 92.360 70.230 ;
        RECT 90.110 69.145 90.440 69.600 ;
        RECT 92.050 69.455 92.370 69.835 ;
        RECT 96.110 69.820 96.410 80.130 ;
        RECT 95.445 69.520 96.410 69.820 ;
        RECT 88.430 68.845 90.440 69.145 ;
        RECT 85.945 67.450 86.275 67.800 ;
        RECT 86.720 67.450 87.050 67.800 ;
        RECT 87.355 67.450 87.685 67.800 ;
        RECT 88.430 67.575 88.730 68.845 ;
        RECT 90.110 68.795 90.440 68.845 ;
        RECT 90.740 68.485 91.060 68.865 ;
        RECT 90.740 68.390 91.050 68.485 ;
        RECT 85.960 66.300 86.260 67.450 ;
        RECT 85.950 65.920 86.270 66.300 ;
        RECT 73.285 58.950 73.615 59.700 ;
        RECT 74.120 59.350 74.450 60.105 ;
        RECT 75.435 59.915 75.765 60.265 ;
        RECT 76.065 59.915 76.395 60.265 ;
        RECT 76.695 59.915 77.025 60.265 ;
        RECT 72.030 57.090 72.345 57.505 ;
        RECT 70.730 56.740 71.060 57.090 ;
        RECT 72.030 56.740 72.360 57.090 ;
        RECT 73.285 56.900 73.615 57.660 ;
        RECT 74.120 57.385 74.450 58.135 ;
        RECT 67.960 51.415 68.290 52.165 ;
        RECT 68.785 51.815 69.115 52.570 ;
        RECT 67.960 49.365 68.290 50.125 ;
        RECT 68.785 49.850 69.115 50.600 ;
        RECT 67.965 47.920 68.295 48.670 ;
        RECT 68.785 48.550 69.115 49.300 ;
        RECT 67.960 45.165 68.290 45.915 ;
        RECT 68.790 45.815 69.120 46.565 ;
        RECT 67.960 43.880 68.290 44.630 ;
        RECT 68.785 44.280 69.115 45.035 ;
        RECT 62.625 36.345 62.955 37.095 ;
        RECT 63.460 36.745 63.790 37.500 ;
        RECT 64.105 37.310 64.435 37.660 ;
        RECT 62.625 34.295 62.955 35.055 ;
        RECT 63.460 34.780 63.790 35.530 ;
        RECT 62.630 32.850 62.960 33.600 ;
        RECT 63.460 33.480 63.790 34.230 ;
        RECT 62.625 30.095 62.955 30.845 ;
        RECT 63.465 30.745 63.795 31.495 ;
        RECT 62.625 28.810 62.955 29.560 ;
        RECT 63.460 29.210 63.790 29.965 ;
        RECT 62.625 26.760 62.955 27.520 ;
        RECT 63.460 27.245 63.790 27.995 ;
        RECT 61.985 26.015 62.315 26.365 ;
        RECT 62.630 25.315 62.960 26.065 ;
        RECT 63.460 25.945 63.790 26.695 ;
        RECT 61.370 24.490 62.310 24.790 ;
        RECT 60.740 23.655 61.675 23.955 ;
        RECT 57.300 21.275 57.630 22.025 ;
        RECT 58.125 21.675 58.455 22.430 ;
        RECT 59.440 22.240 59.770 22.590 ;
        RECT 60.700 22.240 61.030 22.590 ;
        RECT 56.670 19.065 57.000 19.415 ;
        RECT 57.300 19.225 57.630 19.985 ;
        RECT 58.125 19.710 58.455 20.460 ;
        RECT 57.305 17.780 57.635 18.530 ;
        RECT 58.125 18.410 58.455 19.160 ;
        RECT 57.300 15.025 57.630 15.775 ;
        RECT 58.130 15.675 58.460 16.425 ;
        RECT 59.455 15.055 59.755 22.240 ;
        RECT 60.715 19.420 61.015 22.240 ;
        RECT 60.070 19.065 60.400 19.415 ;
        RECT 60.700 19.070 61.030 19.420 ;
        RECT 60.085 15.055 60.385 19.065 ;
        RECT 60.715 15.055 61.015 19.070 ;
        RECT 57.300 13.740 57.630 14.490 ;
        RECT 58.125 14.140 58.455 14.895 ;
        RECT 59.440 14.705 59.770 15.055 ;
        RECT 60.070 14.705 60.400 15.055 ;
        RECT 60.700 14.705 61.030 15.055 ;
        RECT 55.400 9.750 55.700 11.535 ;
        RECT 56.035 11.530 56.365 11.880 ;
        RECT 57.300 11.620 57.630 12.450 ;
        RECT 58.125 12.175 58.455 12.925 ;
        RECT 60.085 11.880 60.385 14.705 ;
        RECT 56.680 11.310 57.630 11.620 ;
        RECT 56.680 10.610 56.990 11.310 ;
        RECT 56.670 10.240 57.000 10.610 ;
        RECT 57.305 10.245 57.635 10.995 ;
        RECT 58.125 10.875 58.455 11.625 ;
        RECT 60.070 11.530 60.400 11.880 ;
        RECT 60.710 11.535 61.040 11.885 ;
        RECT 61.375 11.880 61.675 23.655 ;
        RECT 62.010 19.415 62.310 24.490 ;
        RECT 62.625 22.560 62.955 23.310 ;
        RECT 63.465 23.210 63.795 23.960 ;
        RECT 64.120 23.090 64.420 37.310 ;
        RECT 64.795 37.155 65.095 37.795 ;
        RECT 65.420 37.660 65.720 38.075 ;
        RECT 66.075 37.660 66.375 41.675 ;
        RECT 67.320 41.670 67.650 42.020 ;
        RECT 67.960 41.830 68.290 42.590 ;
        RECT 68.785 42.315 69.115 43.065 ;
        RECT 65.405 37.310 66.375 37.660 ;
        RECT 64.780 36.805 65.110 37.155 ;
        RECT 64.795 35.125 65.095 36.805 ;
        RECT 64.780 34.775 65.110 35.125 ;
        RECT 64.795 30.835 65.095 34.775 ;
        RECT 65.405 34.135 65.735 34.485 ;
        RECT 64.780 30.485 65.110 30.835 ;
        RECT 65.420 30.125 65.720 34.135 ;
        RECT 64.775 29.775 65.105 30.125 ;
        RECT 65.405 29.775 65.735 30.125 ;
        RECT 64.105 22.740 64.435 23.090 ;
        RECT 64.790 22.590 65.090 29.775 ;
        RECT 65.420 26.950 65.720 29.775 ;
        RECT 65.405 26.600 65.735 26.950 ;
        RECT 66.075 23.955 66.375 37.310 ;
        RECT 66.690 34.135 67.020 34.485 ;
        RECT 66.705 27.365 67.005 34.135 ;
        RECT 66.705 26.950 67.020 27.365 ;
        RECT 66.705 26.600 67.035 26.950 ;
        RECT 66.705 24.790 67.005 26.600 ;
        RECT 67.335 26.365 67.635 41.670 ;
        RECT 67.965 40.385 68.295 41.135 ;
        RECT 68.785 41.015 69.115 41.765 ;
        RECT 67.960 37.630 68.290 38.380 ;
        RECT 68.790 38.280 69.120 39.030 ;
        RECT 69.445 37.660 69.745 52.960 ;
        RECT 70.115 52.730 70.430 53.145 ;
        RECT 70.115 52.380 70.445 52.730 ;
        RECT 71.360 52.380 71.690 52.730 ;
        RECT 70.115 45.195 70.415 52.380 ;
        RECT 71.375 49.560 71.675 52.380 ;
        RECT 70.730 49.205 71.060 49.555 ;
        RECT 71.360 49.210 71.690 49.560 ;
        RECT 72.030 49.555 72.330 56.740 ;
        RECT 72.645 56.235 72.975 56.585 ;
        RECT 70.745 45.195 71.045 49.205 ;
        RECT 71.375 45.195 71.675 49.210 ;
        RECT 72.015 49.205 72.345 49.555 ;
        RECT 70.100 44.845 70.430 45.195 ;
        RECT 70.730 44.845 71.060 45.195 ;
        RECT 71.360 44.845 71.690 45.195 ;
        RECT 70.745 42.020 71.045 44.845 ;
        RECT 70.730 41.670 71.060 42.020 ;
        RECT 71.385 41.675 71.715 42.025 ;
        RECT 72.660 42.020 72.960 56.235 ;
        RECT 73.290 55.455 73.620 56.205 ;
        RECT 74.120 56.085 74.450 56.835 ;
        RECT 73.285 52.700 73.615 53.450 ;
        RECT 74.125 53.350 74.455 54.100 ;
        RECT 74.765 52.960 75.095 53.310 ;
        RECT 75.450 53.145 75.750 59.915 ;
        RECT 76.080 57.090 76.380 59.915 ;
        RECT 77.365 57.505 77.665 64.275 ;
        RECT 78.625 62.990 78.955 63.740 ;
        RECT 79.445 63.620 79.775 64.370 ;
        RECT 81.390 64.275 81.720 64.625 ;
        RECT 82.020 64.280 82.350 64.630 ;
        RECT 78.620 60.235 78.950 60.985 ;
        RECT 79.450 60.885 79.780 61.635 ;
        RECT 81.405 60.265 81.705 64.275 ;
        RECT 82.035 60.265 82.335 64.280 ;
        RECT 82.675 64.275 83.005 64.625 ;
        RECT 83.945 64.435 84.275 65.195 ;
        RECT 84.780 64.920 85.110 65.670 ;
        RECT 87.370 64.630 87.670 67.450 ;
        RECT 88.420 67.195 88.740 67.575 ;
        RECT 89.280 67.535 89.610 68.270 ;
        RECT 90.105 68.090 91.050 68.390 ;
        RECT 89.280 66.485 89.610 67.235 ;
        RECT 90.105 66.935 90.435 68.090 ;
        RECT 92.060 67.800 92.360 69.455 ;
        RECT 95.445 68.795 95.775 69.520 ;
        RECT 96.740 68.495 97.040 80.515 ;
        RECT 106.770 79.720 107.070 80.135 ;
        RECT 107.400 80.090 107.700 80.505 ;
        RECT 107.385 79.740 107.715 80.090 ;
        RECT 106.755 79.370 107.085 79.720 ;
        RECT 97.385 73.385 97.705 73.765 ;
        RECT 91.270 67.450 91.600 67.800 ;
        RECT 92.045 67.450 92.375 67.800 ;
        RECT 92.680 67.450 93.010 67.800 ;
        RECT 94.605 67.535 94.935 68.270 ;
        RECT 95.440 68.195 97.040 68.495 ;
        RECT 91.285 66.300 91.585 67.450 ;
        RECT 91.275 65.920 91.595 66.300 ;
        RECT 78.620 58.950 78.950 59.700 ;
        RECT 79.445 59.350 79.775 60.105 ;
        RECT 80.760 59.915 81.090 60.265 ;
        RECT 81.390 59.915 81.720 60.265 ;
        RECT 82.020 59.915 82.350 60.265 ;
        RECT 77.365 57.090 77.680 57.505 ;
        RECT 76.065 56.740 76.395 57.090 ;
        RECT 77.365 56.740 77.695 57.090 ;
        RECT 78.620 56.900 78.950 57.660 ;
        RECT 79.445 57.385 79.775 58.135 ;
        RECT 73.285 51.415 73.615 52.165 ;
        RECT 74.120 51.815 74.450 52.570 ;
        RECT 73.285 49.365 73.615 50.125 ;
        RECT 74.120 49.850 74.450 50.600 ;
        RECT 73.290 47.920 73.620 48.670 ;
        RECT 74.120 48.550 74.450 49.300 ;
        RECT 73.285 45.165 73.615 45.915 ;
        RECT 74.125 45.815 74.455 46.565 ;
        RECT 73.285 43.880 73.615 44.630 ;
        RECT 74.120 44.280 74.450 45.035 ;
        RECT 67.960 36.345 68.290 37.095 ;
        RECT 68.785 36.745 69.115 37.500 ;
        RECT 69.430 37.310 69.760 37.660 ;
        RECT 67.960 34.295 68.290 35.055 ;
        RECT 68.785 34.780 69.115 35.530 ;
        RECT 67.965 32.850 68.295 33.600 ;
        RECT 68.785 33.480 69.115 34.230 ;
        RECT 67.960 30.095 68.290 30.845 ;
        RECT 68.790 30.745 69.120 31.495 ;
        RECT 67.960 28.810 68.290 29.560 ;
        RECT 68.785 29.210 69.115 29.965 ;
        RECT 67.960 26.760 68.290 27.520 ;
        RECT 68.785 27.245 69.115 27.995 ;
        RECT 67.320 26.015 67.650 26.365 ;
        RECT 67.965 25.315 68.295 26.065 ;
        RECT 68.785 25.945 69.115 26.695 ;
        RECT 66.705 24.490 67.645 24.790 ;
        RECT 66.075 23.655 67.010 23.955 ;
        RECT 62.625 21.275 62.955 22.025 ;
        RECT 63.460 21.675 63.790 22.430 ;
        RECT 64.775 22.240 65.105 22.590 ;
        RECT 66.035 22.240 66.365 22.590 ;
        RECT 61.995 19.065 62.325 19.415 ;
        RECT 62.625 19.225 62.955 19.985 ;
        RECT 63.460 19.710 63.790 20.460 ;
        RECT 62.630 17.780 62.960 18.530 ;
        RECT 63.460 18.410 63.790 19.160 ;
        RECT 62.625 15.025 62.955 15.775 ;
        RECT 63.465 15.675 63.795 16.425 ;
        RECT 64.790 15.055 65.090 22.240 ;
        RECT 66.050 19.420 66.350 22.240 ;
        RECT 65.405 19.065 65.735 19.415 ;
        RECT 66.035 19.070 66.365 19.420 ;
        RECT 65.420 15.055 65.720 19.065 ;
        RECT 66.050 15.055 66.350 19.070 ;
        RECT 62.625 13.740 62.955 14.490 ;
        RECT 63.460 14.140 63.790 14.895 ;
        RECT 64.775 14.705 65.105 15.055 ;
        RECT 65.405 14.705 65.735 15.055 ;
        RECT 66.035 14.705 66.365 15.055 ;
        RECT 50.055 9.210 50.375 9.590 ;
        RECT 55.390 9.370 55.710 9.750 ;
        RECT 60.725 9.590 61.025 11.535 ;
        RECT 61.360 11.530 61.690 11.880 ;
        RECT 62.625 11.690 62.955 12.450 ;
        RECT 63.460 12.175 63.790 12.925 ;
        RECT 65.420 11.880 65.720 14.705 ;
        RECT 62.630 10.245 62.960 10.995 ;
        RECT 63.460 10.875 63.790 11.625 ;
        RECT 65.405 11.530 65.735 11.880 ;
        RECT 66.045 11.535 66.375 11.885 ;
        RECT 66.710 11.880 67.010 23.655 ;
        RECT 67.345 19.415 67.645 24.490 ;
        RECT 67.960 22.560 68.290 23.310 ;
        RECT 68.790 23.210 69.120 23.960 ;
        RECT 69.445 23.090 69.745 37.310 ;
        RECT 70.120 37.155 70.420 37.795 ;
        RECT 70.745 37.660 71.045 38.075 ;
        RECT 71.400 37.660 71.700 41.675 ;
        RECT 72.645 41.670 72.975 42.020 ;
        RECT 73.285 41.830 73.615 42.590 ;
        RECT 74.120 42.315 74.450 43.065 ;
        RECT 70.730 37.310 71.700 37.660 ;
        RECT 70.105 36.805 70.435 37.155 ;
        RECT 70.120 35.125 70.420 36.805 ;
        RECT 70.105 34.775 70.435 35.125 ;
        RECT 70.120 30.835 70.420 34.775 ;
        RECT 70.730 34.135 71.060 34.485 ;
        RECT 70.105 30.485 70.435 30.835 ;
        RECT 70.745 30.125 71.045 34.135 ;
        RECT 70.100 29.775 70.430 30.125 ;
        RECT 70.730 29.775 71.060 30.125 ;
        RECT 69.430 22.740 69.760 23.090 ;
        RECT 70.115 22.590 70.415 29.775 ;
        RECT 70.745 26.950 71.045 29.775 ;
        RECT 70.730 26.600 71.060 26.950 ;
        RECT 71.400 23.955 71.700 37.310 ;
        RECT 72.015 34.135 72.345 34.485 ;
        RECT 72.030 27.365 72.330 34.135 ;
        RECT 72.030 26.950 72.345 27.365 ;
        RECT 72.030 26.600 72.360 26.950 ;
        RECT 72.030 24.790 72.330 26.600 ;
        RECT 72.660 26.365 72.960 41.670 ;
        RECT 73.290 40.385 73.620 41.135 ;
        RECT 74.120 41.015 74.450 41.765 ;
        RECT 73.285 37.630 73.615 38.380 ;
        RECT 74.125 38.280 74.455 39.030 ;
        RECT 74.780 37.660 75.080 52.960 ;
        RECT 75.450 52.730 75.765 53.145 ;
        RECT 75.450 52.380 75.780 52.730 ;
        RECT 76.695 52.380 77.025 52.730 ;
        RECT 75.450 45.195 75.750 52.380 ;
        RECT 76.710 49.560 77.010 52.380 ;
        RECT 76.065 49.205 76.395 49.555 ;
        RECT 76.695 49.210 77.025 49.560 ;
        RECT 77.365 49.555 77.665 56.740 ;
        RECT 77.980 56.235 78.310 56.585 ;
        RECT 76.080 45.195 76.380 49.205 ;
        RECT 76.710 45.195 77.010 49.210 ;
        RECT 77.350 49.205 77.680 49.555 ;
        RECT 75.435 44.845 75.765 45.195 ;
        RECT 76.065 44.845 76.395 45.195 ;
        RECT 76.695 44.845 77.025 45.195 ;
        RECT 76.080 42.020 76.380 44.845 ;
        RECT 76.065 41.670 76.395 42.020 ;
        RECT 76.720 41.675 77.050 42.025 ;
        RECT 77.995 42.020 78.295 56.235 ;
        RECT 78.625 55.455 78.955 56.205 ;
        RECT 79.445 56.085 79.775 56.835 ;
        RECT 78.620 52.700 78.950 53.450 ;
        RECT 79.450 53.350 79.780 54.100 ;
        RECT 80.090 52.960 80.420 53.310 ;
        RECT 80.775 53.145 81.075 59.915 ;
        RECT 81.405 57.090 81.705 59.915 ;
        RECT 82.690 57.505 82.990 64.275 ;
        RECT 83.950 62.990 84.280 63.740 ;
        RECT 84.780 63.620 85.110 64.370 ;
        RECT 86.725 64.275 87.055 64.625 ;
        RECT 87.355 64.280 87.685 64.630 ;
        RECT 83.945 60.235 84.275 60.985 ;
        RECT 84.785 60.885 85.115 61.635 ;
        RECT 86.740 60.265 87.040 64.275 ;
        RECT 87.370 60.265 87.670 64.280 ;
        RECT 88.010 64.275 88.340 64.625 ;
        RECT 89.280 64.435 89.610 65.195 ;
        RECT 90.105 64.920 90.435 65.670 ;
        RECT 92.695 64.630 92.995 67.450 ;
        RECT 94.605 66.485 94.935 67.235 ;
        RECT 95.440 66.935 95.770 68.195 ;
        RECT 97.395 67.800 97.695 73.385 ;
        RECT 102.720 69.835 103.020 70.230 ;
        RECT 100.770 68.795 101.100 69.600 ;
        RECT 102.710 69.455 103.030 69.835 ;
        RECT 106.770 69.820 107.070 79.370 ;
        RECT 106.105 69.520 107.070 69.820 ;
        RECT 100.770 68.485 101.090 68.795 ;
        RECT 97.380 67.450 97.710 67.800 ;
        RECT 98.015 67.450 98.345 67.800 ;
        RECT 99.940 67.535 100.270 68.270 ;
        RECT 100.780 67.670 101.080 67.970 ;
        RECT 102.720 67.800 103.020 69.455 ;
        RECT 106.105 68.795 106.435 69.520 ;
        RECT 107.400 68.495 107.700 79.740 ;
        RECT 108.045 73.385 108.365 73.765 ;
        RECT 83.945 58.950 84.275 59.700 ;
        RECT 84.780 59.350 85.110 60.105 ;
        RECT 86.095 59.915 86.425 60.265 ;
        RECT 86.725 59.915 87.055 60.265 ;
        RECT 87.355 59.915 87.685 60.265 ;
        RECT 82.690 57.090 83.005 57.505 ;
        RECT 81.390 56.740 81.720 57.090 ;
        RECT 82.690 56.740 83.020 57.090 ;
        RECT 83.945 56.900 84.275 57.660 ;
        RECT 84.780 57.385 85.110 58.135 ;
        RECT 78.620 51.415 78.950 52.165 ;
        RECT 79.445 51.815 79.775 52.570 ;
        RECT 78.620 49.365 78.950 50.125 ;
        RECT 79.445 49.850 79.775 50.600 ;
        RECT 78.625 47.920 78.955 48.670 ;
        RECT 79.445 48.550 79.775 49.300 ;
        RECT 78.620 45.165 78.950 45.915 ;
        RECT 79.450 45.815 79.780 46.565 ;
        RECT 78.620 43.880 78.950 44.630 ;
        RECT 79.445 44.280 79.775 45.035 ;
        RECT 73.285 36.345 73.615 37.095 ;
        RECT 74.120 36.745 74.450 37.500 ;
        RECT 74.765 37.310 75.095 37.660 ;
        RECT 73.285 34.295 73.615 35.055 ;
        RECT 74.120 34.780 74.450 35.530 ;
        RECT 73.290 32.850 73.620 33.600 ;
        RECT 74.120 33.480 74.450 34.230 ;
        RECT 73.285 30.095 73.615 30.845 ;
        RECT 74.125 30.745 74.455 31.495 ;
        RECT 73.285 28.810 73.615 29.560 ;
        RECT 74.120 29.210 74.450 29.965 ;
        RECT 73.285 26.760 73.615 27.520 ;
        RECT 74.120 27.245 74.450 27.995 ;
        RECT 72.645 26.015 72.975 26.365 ;
        RECT 73.290 25.315 73.620 26.065 ;
        RECT 74.120 25.945 74.450 26.695 ;
        RECT 72.030 24.490 72.970 24.790 ;
        RECT 71.400 23.655 72.335 23.955 ;
        RECT 67.960 21.275 68.290 22.025 ;
        RECT 68.785 21.675 69.115 22.430 ;
        RECT 70.100 22.240 70.430 22.590 ;
        RECT 71.360 22.240 71.690 22.590 ;
        RECT 67.330 19.065 67.660 19.415 ;
        RECT 67.960 19.225 68.290 19.985 ;
        RECT 68.785 19.710 69.115 20.460 ;
        RECT 67.965 17.780 68.295 18.530 ;
        RECT 68.785 18.410 69.115 19.160 ;
        RECT 67.960 15.025 68.290 15.775 ;
        RECT 68.790 15.675 69.120 16.425 ;
        RECT 70.115 15.055 70.415 22.240 ;
        RECT 71.375 19.420 71.675 22.240 ;
        RECT 70.730 19.065 71.060 19.415 ;
        RECT 71.360 19.070 71.690 19.420 ;
        RECT 70.745 15.055 71.045 19.065 ;
        RECT 71.375 15.055 71.675 19.070 ;
        RECT 67.960 13.740 68.290 14.490 ;
        RECT 68.785 14.140 69.115 14.895 ;
        RECT 70.100 14.705 70.430 15.055 ;
        RECT 70.730 14.705 71.060 15.055 ;
        RECT 71.360 14.705 71.690 15.055 ;
        RECT 66.060 9.750 66.360 11.535 ;
        RECT 66.695 11.530 67.025 11.880 ;
        RECT 67.960 11.620 68.290 12.450 ;
        RECT 68.785 12.175 69.115 12.925 ;
        RECT 70.745 11.880 71.045 14.705 ;
        RECT 67.340 11.310 68.290 11.620 ;
        RECT 67.340 10.610 67.650 11.310 ;
        RECT 67.330 10.240 67.660 10.610 ;
        RECT 67.965 10.245 68.295 10.995 ;
        RECT 68.785 10.875 69.115 11.625 ;
        RECT 70.730 11.530 71.060 11.880 ;
        RECT 71.370 11.535 71.700 11.885 ;
        RECT 72.035 11.880 72.335 23.655 ;
        RECT 72.670 19.415 72.970 24.490 ;
        RECT 73.285 22.560 73.615 23.310 ;
        RECT 74.125 23.210 74.455 23.960 ;
        RECT 74.780 23.090 75.080 37.310 ;
        RECT 75.455 37.155 75.755 37.795 ;
        RECT 76.080 37.660 76.380 38.075 ;
        RECT 76.735 37.660 77.035 41.675 ;
        RECT 77.980 41.670 78.310 42.020 ;
        RECT 78.620 41.830 78.950 42.590 ;
        RECT 79.445 42.315 79.775 43.065 ;
        RECT 76.065 37.310 77.035 37.660 ;
        RECT 75.440 36.805 75.770 37.155 ;
        RECT 75.455 35.125 75.755 36.805 ;
        RECT 75.440 34.775 75.770 35.125 ;
        RECT 75.455 30.835 75.755 34.775 ;
        RECT 76.065 34.135 76.395 34.485 ;
        RECT 75.440 30.485 75.770 30.835 ;
        RECT 76.080 30.125 76.380 34.135 ;
        RECT 75.435 29.775 75.765 30.125 ;
        RECT 76.065 29.775 76.395 30.125 ;
        RECT 74.765 22.740 75.095 23.090 ;
        RECT 75.450 22.590 75.750 29.775 ;
        RECT 76.080 26.950 76.380 29.775 ;
        RECT 76.065 26.600 76.395 26.950 ;
        RECT 76.735 23.955 77.035 37.310 ;
        RECT 77.350 34.135 77.680 34.485 ;
        RECT 77.365 27.365 77.665 34.135 ;
        RECT 77.365 26.950 77.680 27.365 ;
        RECT 77.365 26.600 77.695 26.950 ;
        RECT 77.365 24.790 77.665 26.600 ;
        RECT 77.995 26.365 78.295 41.670 ;
        RECT 78.625 40.385 78.955 41.135 ;
        RECT 79.445 41.015 79.775 41.765 ;
        RECT 78.620 37.630 78.950 38.380 ;
        RECT 79.450 38.280 79.780 39.030 ;
        RECT 80.105 37.660 80.405 52.960 ;
        RECT 80.775 52.730 81.090 53.145 ;
        RECT 80.775 52.380 81.105 52.730 ;
        RECT 82.020 52.380 82.350 52.730 ;
        RECT 80.775 45.195 81.075 52.380 ;
        RECT 82.035 49.560 82.335 52.380 ;
        RECT 81.390 49.205 81.720 49.555 ;
        RECT 82.020 49.210 82.350 49.560 ;
        RECT 82.690 49.555 82.990 56.740 ;
        RECT 83.305 56.235 83.635 56.585 ;
        RECT 81.405 45.195 81.705 49.205 ;
        RECT 82.035 45.195 82.335 49.210 ;
        RECT 82.675 49.205 83.005 49.555 ;
        RECT 80.760 44.845 81.090 45.195 ;
        RECT 81.390 44.845 81.720 45.195 ;
        RECT 82.020 44.845 82.350 45.195 ;
        RECT 81.405 42.020 81.705 44.845 ;
        RECT 81.390 41.670 81.720 42.020 ;
        RECT 82.045 41.675 82.375 42.025 ;
        RECT 83.320 42.020 83.620 56.235 ;
        RECT 83.950 55.455 84.280 56.205 ;
        RECT 84.780 56.085 85.110 56.835 ;
        RECT 83.945 52.700 84.275 53.450 ;
        RECT 84.785 53.350 85.115 54.100 ;
        RECT 85.425 52.960 85.755 53.310 ;
        RECT 86.110 53.145 86.410 59.915 ;
        RECT 86.740 57.090 87.040 59.915 ;
        RECT 88.025 57.505 88.325 64.275 ;
        RECT 89.285 62.990 89.615 63.740 ;
        RECT 90.105 63.620 90.435 64.370 ;
        RECT 92.050 64.275 92.380 64.625 ;
        RECT 92.680 64.280 93.010 64.630 ;
        RECT 89.280 60.235 89.610 60.985 ;
        RECT 90.110 60.885 90.440 61.635 ;
        RECT 92.065 60.265 92.365 64.275 ;
        RECT 92.695 60.265 92.995 64.280 ;
        RECT 93.335 64.275 93.665 64.625 ;
        RECT 94.605 64.435 94.935 65.195 ;
        RECT 95.440 64.920 95.770 65.670 ;
        RECT 98.030 64.630 98.330 67.450 ;
        RECT 99.940 66.485 100.270 67.235 ;
        RECT 100.765 66.935 101.095 67.670 ;
        RECT 101.930 67.450 102.260 67.800 ;
        RECT 102.705 67.450 103.035 67.800 ;
        RECT 103.340 67.450 103.670 67.800 ;
        RECT 105.265 67.535 105.595 68.270 ;
        RECT 106.100 68.195 107.700 68.495 ;
        RECT 101.945 66.300 102.245 67.450 ;
        RECT 101.935 65.920 102.255 66.300 ;
        RECT 89.280 58.950 89.610 59.700 ;
        RECT 90.105 59.350 90.435 60.105 ;
        RECT 91.420 59.915 91.750 60.265 ;
        RECT 92.050 59.915 92.380 60.265 ;
        RECT 92.680 59.915 93.010 60.265 ;
        RECT 88.025 57.090 88.340 57.505 ;
        RECT 86.725 56.740 87.055 57.090 ;
        RECT 88.025 56.740 88.355 57.090 ;
        RECT 89.280 56.900 89.610 57.660 ;
        RECT 90.105 57.385 90.435 58.135 ;
        RECT 83.945 51.415 84.275 52.165 ;
        RECT 84.780 51.815 85.110 52.570 ;
        RECT 83.945 49.365 84.275 50.125 ;
        RECT 84.780 49.850 85.110 50.600 ;
        RECT 83.950 47.920 84.280 48.670 ;
        RECT 84.780 48.550 85.110 49.300 ;
        RECT 83.945 45.165 84.275 45.915 ;
        RECT 84.785 45.815 85.115 46.565 ;
        RECT 83.945 43.880 84.275 44.630 ;
        RECT 84.780 44.280 85.110 45.035 ;
        RECT 78.620 36.345 78.950 37.095 ;
        RECT 79.445 36.745 79.775 37.500 ;
        RECT 80.090 37.310 80.420 37.660 ;
        RECT 78.620 34.295 78.950 35.055 ;
        RECT 79.445 34.780 79.775 35.530 ;
        RECT 78.625 32.850 78.955 33.600 ;
        RECT 79.445 33.480 79.775 34.230 ;
        RECT 78.620 30.095 78.950 30.845 ;
        RECT 79.450 30.745 79.780 31.495 ;
        RECT 78.620 28.810 78.950 29.560 ;
        RECT 79.445 29.210 79.775 29.965 ;
        RECT 78.620 26.760 78.950 27.520 ;
        RECT 79.445 27.245 79.775 27.995 ;
        RECT 77.980 26.015 78.310 26.365 ;
        RECT 78.625 25.315 78.955 26.065 ;
        RECT 79.445 25.945 79.775 26.695 ;
        RECT 77.365 24.490 78.305 24.790 ;
        RECT 76.735 23.655 77.670 23.955 ;
        RECT 73.285 21.275 73.615 22.025 ;
        RECT 74.120 21.675 74.450 22.430 ;
        RECT 75.435 22.240 75.765 22.590 ;
        RECT 76.695 22.240 77.025 22.590 ;
        RECT 72.655 19.065 72.985 19.415 ;
        RECT 73.285 19.225 73.615 19.985 ;
        RECT 74.120 19.710 74.450 20.460 ;
        RECT 73.290 17.780 73.620 18.530 ;
        RECT 74.120 18.410 74.450 19.160 ;
        RECT 73.285 15.025 73.615 15.775 ;
        RECT 74.125 15.675 74.455 16.425 ;
        RECT 75.450 15.055 75.750 22.240 ;
        RECT 76.710 19.420 77.010 22.240 ;
        RECT 76.065 19.065 76.395 19.415 ;
        RECT 76.695 19.070 77.025 19.420 ;
        RECT 76.080 15.055 76.380 19.065 ;
        RECT 76.710 15.055 77.010 19.070 ;
        RECT 73.285 13.740 73.615 14.490 ;
        RECT 74.120 14.140 74.450 14.895 ;
        RECT 75.435 14.705 75.765 15.055 ;
        RECT 76.065 14.705 76.395 15.055 ;
        RECT 76.695 14.705 77.025 15.055 ;
        RECT 60.715 9.210 61.035 9.590 ;
        RECT 66.050 9.370 66.370 9.750 ;
        RECT 71.385 9.590 71.685 11.535 ;
        RECT 72.020 11.530 72.350 11.880 ;
        RECT 73.285 11.690 73.615 12.450 ;
        RECT 74.120 12.175 74.450 12.925 ;
        RECT 76.080 11.880 76.380 14.705 ;
        RECT 73.290 10.245 73.620 10.995 ;
        RECT 74.120 10.875 74.450 11.625 ;
        RECT 76.065 11.530 76.395 11.880 ;
        RECT 76.705 11.535 77.035 11.885 ;
        RECT 77.370 11.880 77.670 23.655 ;
        RECT 78.005 19.415 78.305 24.490 ;
        RECT 78.620 22.560 78.950 23.310 ;
        RECT 79.450 23.210 79.780 23.960 ;
        RECT 80.105 23.090 80.405 37.310 ;
        RECT 80.780 37.155 81.080 37.795 ;
        RECT 81.405 37.660 81.705 38.075 ;
        RECT 82.060 37.660 82.360 41.675 ;
        RECT 83.305 41.670 83.635 42.020 ;
        RECT 83.945 41.830 84.275 42.590 ;
        RECT 84.780 42.315 85.110 43.065 ;
        RECT 81.390 37.310 82.360 37.660 ;
        RECT 80.765 36.805 81.095 37.155 ;
        RECT 80.780 35.125 81.080 36.805 ;
        RECT 80.765 34.775 81.095 35.125 ;
        RECT 80.780 30.835 81.080 34.775 ;
        RECT 81.390 34.135 81.720 34.485 ;
        RECT 80.765 30.485 81.095 30.835 ;
        RECT 81.405 30.125 81.705 34.135 ;
        RECT 80.760 29.775 81.090 30.125 ;
        RECT 81.390 29.775 81.720 30.125 ;
        RECT 80.090 22.740 80.420 23.090 ;
        RECT 80.775 22.590 81.075 29.775 ;
        RECT 81.405 26.950 81.705 29.775 ;
        RECT 81.390 26.600 81.720 26.950 ;
        RECT 82.060 23.955 82.360 37.310 ;
        RECT 82.675 34.135 83.005 34.485 ;
        RECT 82.690 27.365 82.990 34.135 ;
        RECT 82.690 26.950 83.005 27.365 ;
        RECT 82.690 26.600 83.020 26.950 ;
        RECT 82.690 24.790 82.990 26.600 ;
        RECT 83.320 26.365 83.620 41.670 ;
        RECT 83.950 40.385 84.280 41.135 ;
        RECT 84.780 41.015 85.110 41.765 ;
        RECT 83.945 37.630 84.275 38.380 ;
        RECT 84.785 38.280 85.115 39.030 ;
        RECT 85.440 37.660 85.740 52.960 ;
        RECT 86.110 52.730 86.425 53.145 ;
        RECT 86.110 52.380 86.440 52.730 ;
        RECT 87.355 52.380 87.685 52.730 ;
        RECT 86.110 45.195 86.410 52.380 ;
        RECT 87.370 49.560 87.670 52.380 ;
        RECT 86.725 49.205 87.055 49.555 ;
        RECT 87.355 49.210 87.685 49.560 ;
        RECT 88.025 49.555 88.325 56.740 ;
        RECT 88.640 56.235 88.970 56.585 ;
        RECT 86.740 45.195 87.040 49.205 ;
        RECT 87.370 45.195 87.670 49.210 ;
        RECT 88.010 49.205 88.340 49.555 ;
        RECT 86.095 44.845 86.425 45.195 ;
        RECT 86.725 44.845 87.055 45.195 ;
        RECT 87.355 44.845 87.685 45.195 ;
        RECT 86.740 42.020 87.040 44.845 ;
        RECT 86.725 41.670 87.055 42.020 ;
        RECT 87.380 41.675 87.710 42.025 ;
        RECT 88.655 42.020 88.955 56.235 ;
        RECT 89.285 55.455 89.615 56.205 ;
        RECT 90.105 56.085 90.435 56.835 ;
        RECT 89.280 52.700 89.610 53.450 ;
        RECT 90.110 53.350 90.440 54.100 ;
        RECT 90.750 52.960 91.080 53.310 ;
        RECT 91.435 53.145 91.735 59.915 ;
        RECT 92.065 57.090 92.365 59.915 ;
        RECT 93.350 57.505 93.650 64.275 ;
        RECT 94.610 62.990 94.940 63.740 ;
        RECT 95.440 63.620 95.770 64.370 ;
        RECT 97.385 64.275 97.715 64.625 ;
        RECT 98.015 64.280 98.345 64.630 ;
        RECT 94.605 60.235 94.935 60.985 ;
        RECT 95.445 60.885 95.775 61.635 ;
        RECT 97.400 60.265 97.700 64.275 ;
        RECT 98.030 60.265 98.330 64.280 ;
        RECT 98.670 64.275 99.000 64.625 ;
        RECT 99.940 64.435 100.270 65.195 ;
        RECT 100.765 64.920 101.095 65.670 ;
        RECT 103.355 64.630 103.655 67.450 ;
        RECT 105.265 66.485 105.595 67.235 ;
        RECT 106.100 66.935 106.430 68.195 ;
        RECT 108.055 67.800 108.355 73.385 ;
        RECT 113.380 69.835 113.680 70.230 ;
        RECT 111.430 69.145 111.760 69.600 ;
        RECT 113.370 69.455 113.690 69.835 ;
        RECT 109.750 68.845 111.760 69.145 ;
        RECT 107.265 67.450 107.595 67.800 ;
        RECT 108.040 67.450 108.370 67.800 ;
        RECT 108.675 67.450 109.005 67.800 ;
        RECT 109.750 67.575 110.050 68.845 ;
        RECT 111.430 68.795 111.760 68.845 ;
        RECT 112.060 68.485 112.380 68.865 ;
        RECT 112.060 68.390 112.370 68.485 ;
        RECT 107.280 66.300 107.580 67.450 ;
        RECT 107.270 65.920 107.590 66.300 ;
        RECT 94.605 58.950 94.935 59.700 ;
        RECT 95.440 59.350 95.770 60.105 ;
        RECT 96.755 59.915 97.085 60.265 ;
        RECT 97.385 59.915 97.715 60.265 ;
        RECT 98.015 59.915 98.345 60.265 ;
        RECT 93.350 57.090 93.665 57.505 ;
        RECT 92.050 56.740 92.380 57.090 ;
        RECT 93.350 56.740 93.680 57.090 ;
        RECT 94.605 56.900 94.935 57.660 ;
        RECT 95.440 57.385 95.770 58.135 ;
        RECT 89.280 51.415 89.610 52.165 ;
        RECT 90.105 51.815 90.435 52.570 ;
        RECT 89.280 49.365 89.610 50.125 ;
        RECT 90.105 49.850 90.435 50.600 ;
        RECT 89.285 47.920 89.615 48.670 ;
        RECT 90.105 48.550 90.435 49.300 ;
        RECT 89.280 45.165 89.610 45.915 ;
        RECT 90.110 45.815 90.440 46.565 ;
        RECT 89.280 43.880 89.610 44.630 ;
        RECT 90.105 44.280 90.435 45.035 ;
        RECT 83.945 36.345 84.275 37.095 ;
        RECT 84.780 36.745 85.110 37.500 ;
        RECT 85.425 37.310 85.755 37.660 ;
        RECT 83.945 34.295 84.275 35.055 ;
        RECT 84.780 34.780 85.110 35.530 ;
        RECT 83.950 32.850 84.280 33.600 ;
        RECT 84.780 33.480 85.110 34.230 ;
        RECT 83.945 30.095 84.275 30.845 ;
        RECT 84.785 30.745 85.115 31.495 ;
        RECT 83.945 28.810 84.275 29.560 ;
        RECT 84.780 29.210 85.110 29.965 ;
        RECT 83.945 26.760 84.275 27.520 ;
        RECT 84.780 27.245 85.110 27.995 ;
        RECT 83.305 26.015 83.635 26.365 ;
        RECT 83.950 25.315 84.280 26.065 ;
        RECT 84.780 25.945 85.110 26.695 ;
        RECT 82.690 24.490 83.630 24.790 ;
        RECT 82.060 23.655 82.995 23.955 ;
        RECT 78.620 21.275 78.950 22.025 ;
        RECT 79.445 21.675 79.775 22.430 ;
        RECT 80.760 22.240 81.090 22.590 ;
        RECT 82.020 22.240 82.350 22.590 ;
        RECT 77.990 19.065 78.320 19.415 ;
        RECT 78.620 19.225 78.950 19.985 ;
        RECT 79.445 19.710 79.775 20.460 ;
        RECT 78.625 17.780 78.955 18.530 ;
        RECT 79.445 18.410 79.775 19.160 ;
        RECT 78.620 15.025 78.950 15.775 ;
        RECT 79.450 15.675 79.780 16.425 ;
        RECT 80.775 15.055 81.075 22.240 ;
        RECT 82.035 19.420 82.335 22.240 ;
        RECT 81.390 19.065 81.720 19.415 ;
        RECT 82.020 19.070 82.350 19.420 ;
        RECT 81.405 15.055 81.705 19.065 ;
        RECT 82.035 15.055 82.335 19.070 ;
        RECT 78.620 13.740 78.950 14.490 ;
        RECT 79.445 14.140 79.775 14.895 ;
        RECT 80.760 14.705 81.090 15.055 ;
        RECT 81.390 14.705 81.720 15.055 ;
        RECT 82.020 14.705 82.350 15.055 ;
        RECT 76.720 9.750 77.020 11.535 ;
        RECT 77.355 11.530 77.685 11.880 ;
        RECT 78.620 11.620 78.950 12.450 ;
        RECT 79.445 12.175 79.775 12.925 ;
        RECT 81.405 11.880 81.705 14.705 ;
        RECT 78.000 11.310 78.950 11.620 ;
        RECT 78.000 10.610 78.310 11.310 ;
        RECT 77.990 10.240 78.320 10.610 ;
        RECT 78.625 10.245 78.955 10.995 ;
        RECT 79.445 10.875 79.775 11.625 ;
        RECT 81.390 11.530 81.720 11.880 ;
        RECT 82.030 11.535 82.360 11.885 ;
        RECT 82.695 11.880 82.995 23.655 ;
        RECT 83.330 19.415 83.630 24.490 ;
        RECT 83.945 22.560 84.275 23.310 ;
        RECT 84.785 23.210 85.115 23.960 ;
        RECT 85.440 23.090 85.740 37.310 ;
        RECT 86.115 37.155 86.415 37.795 ;
        RECT 86.740 37.660 87.040 38.075 ;
        RECT 87.395 37.660 87.695 41.675 ;
        RECT 88.640 41.670 88.970 42.020 ;
        RECT 89.280 41.830 89.610 42.590 ;
        RECT 90.105 42.315 90.435 43.065 ;
        RECT 86.725 37.310 87.695 37.660 ;
        RECT 86.100 36.805 86.430 37.155 ;
        RECT 86.115 35.125 86.415 36.805 ;
        RECT 86.100 34.775 86.430 35.125 ;
        RECT 86.115 30.835 86.415 34.775 ;
        RECT 86.725 34.135 87.055 34.485 ;
        RECT 86.100 30.485 86.430 30.835 ;
        RECT 86.740 30.125 87.040 34.135 ;
        RECT 86.095 29.775 86.425 30.125 ;
        RECT 86.725 29.775 87.055 30.125 ;
        RECT 85.425 22.740 85.755 23.090 ;
        RECT 86.110 22.590 86.410 29.775 ;
        RECT 86.740 26.950 87.040 29.775 ;
        RECT 86.725 26.600 87.055 26.950 ;
        RECT 87.395 23.955 87.695 37.310 ;
        RECT 88.010 34.135 88.340 34.485 ;
        RECT 88.025 27.365 88.325 34.135 ;
        RECT 88.025 26.950 88.340 27.365 ;
        RECT 88.025 26.600 88.355 26.950 ;
        RECT 88.025 24.790 88.325 26.600 ;
        RECT 88.655 26.365 88.955 41.670 ;
        RECT 89.285 40.385 89.615 41.135 ;
        RECT 90.105 41.015 90.435 41.765 ;
        RECT 89.280 37.630 89.610 38.380 ;
        RECT 90.110 38.280 90.440 39.030 ;
        RECT 90.765 37.660 91.065 52.960 ;
        RECT 91.435 52.730 91.750 53.145 ;
        RECT 91.435 52.380 91.765 52.730 ;
        RECT 92.680 52.380 93.010 52.730 ;
        RECT 91.435 45.195 91.735 52.380 ;
        RECT 92.695 49.560 92.995 52.380 ;
        RECT 92.050 49.205 92.380 49.555 ;
        RECT 92.680 49.210 93.010 49.560 ;
        RECT 93.350 49.555 93.650 56.740 ;
        RECT 93.965 56.235 94.295 56.585 ;
        RECT 92.065 45.195 92.365 49.205 ;
        RECT 92.695 45.195 92.995 49.210 ;
        RECT 93.335 49.205 93.665 49.555 ;
        RECT 91.420 44.845 91.750 45.195 ;
        RECT 92.050 44.845 92.380 45.195 ;
        RECT 92.680 44.845 93.010 45.195 ;
        RECT 92.065 42.020 92.365 44.845 ;
        RECT 92.050 41.670 92.380 42.020 ;
        RECT 92.705 41.675 93.035 42.025 ;
        RECT 93.980 42.020 94.280 56.235 ;
        RECT 94.610 55.455 94.940 56.205 ;
        RECT 95.440 56.085 95.770 56.835 ;
        RECT 94.605 52.700 94.935 53.450 ;
        RECT 95.445 53.350 95.775 54.100 ;
        RECT 96.085 52.960 96.415 53.310 ;
        RECT 96.770 53.145 97.070 59.915 ;
        RECT 97.400 57.090 97.700 59.915 ;
        RECT 98.685 57.505 98.985 64.275 ;
        RECT 99.945 62.990 100.275 63.740 ;
        RECT 100.765 63.620 101.095 64.370 ;
        RECT 102.710 64.275 103.040 64.625 ;
        RECT 103.340 64.280 103.670 64.630 ;
        RECT 99.940 60.235 100.270 60.985 ;
        RECT 100.770 60.885 101.100 61.635 ;
        RECT 102.725 60.265 103.025 64.275 ;
        RECT 103.355 60.265 103.655 64.280 ;
        RECT 103.995 64.275 104.325 64.625 ;
        RECT 105.265 64.435 105.595 65.195 ;
        RECT 106.100 64.920 106.430 65.670 ;
        RECT 108.690 64.630 108.990 67.450 ;
        RECT 109.740 67.195 110.060 67.575 ;
        RECT 110.600 67.535 110.930 68.270 ;
        RECT 111.425 68.090 112.370 68.390 ;
        RECT 110.600 66.485 110.930 67.235 ;
        RECT 111.425 66.935 111.755 68.090 ;
        RECT 113.380 67.800 113.680 69.455 ;
        RECT 112.590 67.450 112.920 67.800 ;
        RECT 113.365 67.450 113.695 67.800 ;
        RECT 114.000 67.450 114.330 67.800 ;
        RECT 115.925 67.535 116.255 68.270 ;
        RECT 118.715 67.800 119.015 70.185 ;
        RECT 117.925 67.450 118.255 67.800 ;
        RECT 118.700 67.450 119.030 67.800 ;
        RECT 119.335 67.450 119.665 67.800 ;
        RECT 121.260 67.535 121.590 68.270 ;
        RECT 112.605 66.300 112.905 67.450 ;
        RECT 112.595 65.920 112.915 66.300 ;
        RECT 99.940 58.950 100.270 59.700 ;
        RECT 100.765 59.350 101.095 60.105 ;
        RECT 102.080 59.915 102.410 60.265 ;
        RECT 102.710 59.915 103.040 60.265 ;
        RECT 103.340 59.915 103.670 60.265 ;
        RECT 98.685 57.090 99.000 57.505 ;
        RECT 97.385 56.740 97.715 57.090 ;
        RECT 98.685 56.740 99.015 57.090 ;
        RECT 99.940 56.900 100.270 57.660 ;
        RECT 100.765 57.385 101.095 58.135 ;
        RECT 94.605 51.415 94.935 52.165 ;
        RECT 95.440 51.815 95.770 52.570 ;
        RECT 94.605 49.365 94.935 50.125 ;
        RECT 95.440 49.850 95.770 50.600 ;
        RECT 94.610 47.920 94.940 48.670 ;
        RECT 95.440 48.550 95.770 49.300 ;
        RECT 94.605 45.165 94.935 45.915 ;
        RECT 95.445 45.815 95.775 46.565 ;
        RECT 94.605 43.880 94.935 44.630 ;
        RECT 95.440 44.280 95.770 45.035 ;
        RECT 89.280 36.345 89.610 37.095 ;
        RECT 90.105 36.745 90.435 37.500 ;
        RECT 90.750 37.310 91.080 37.660 ;
        RECT 89.280 34.295 89.610 35.055 ;
        RECT 90.105 34.780 90.435 35.530 ;
        RECT 89.285 32.850 89.615 33.600 ;
        RECT 90.105 33.480 90.435 34.230 ;
        RECT 89.280 30.095 89.610 30.845 ;
        RECT 90.110 30.745 90.440 31.495 ;
        RECT 89.280 28.810 89.610 29.560 ;
        RECT 90.105 29.210 90.435 29.965 ;
        RECT 89.280 26.760 89.610 27.520 ;
        RECT 90.105 27.245 90.435 27.995 ;
        RECT 88.640 26.015 88.970 26.365 ;
        RECT 89.285 25.315 89.615 26.065 ;
        RECT 90.105 25.945 90.435 26.695 ;
        RECT 88.025 24.490 88.965 24.790 ;
        RECT 87.395 23.655 88.330 23.955 ;
        RECT 83.945 21.275 84.275 22.025 ;
        RECT 84.780 21.675 85.110 22.430 ;
        RECT 86.095 22.240 86.425 22.590 ;
        RECT 87.355 22.240 87.685 22.590 ;
        RECT 83.315 19.065 83.645 19.415 ;
        RECT 83.945 19.225 84.275 19.985 ;
        RECT 84.780 19.710 85.110 20.460 ;
        RECT 83.950 17.780 84.280 18.530 ;
        RECT 84.780 18.410 85.110 19.160 ;
        RECT 83.945 15.025 84.275 15.775 ;
        RECT 84.785 15.675 85.115 16.425 ;
        RECT 86.110 15.055 86.410 22.240 ;
        RECT 87.370 19.420 87.670 22.240 ;
        RECT 86.725 19.065 87.055 19.415 ;
        RECT 87.355 19.070 87.685 19.420 ;
        RECT 86.740 15.055 87.040 19.065 ;
        RECT 87.370 15.055 87.670 19.070 ;
        RECT 83.945 13.740 84.275 14.490 ;
        RECT 84.780 14.140 85.110 14.895 ;
        RECT 86.095 14.705 86.425 15.055 ;
        RECT 86.725 14.705 87.055 15.055 ;
        RECT 87.355 14.705 87.685 15.055 ;
        RECT 71.375 9.210 71.695 9.590 ;
        RECT 76.710 9.370 77.030 9.750 ;
        RECT 82.045 9.590 82.345 11.535 ;
        RECT 82.680 11.530 83.010 11.880 ;
        RECT 83.945 11.690 84.275 12.450 ;
        RECT 84.780 12.175 85.110 12.925 ;
        RECT 86.740 11.880 87.040 14.705 ;
        RECT 83.950 10.245 84.280 10.995 ;
        RECT 84.780 10.875 85.110 11.625 ;
        RECT 86.725 11.530 87.055 11.880 ;
        RECT 87.365 11.535 87.695 11.885 ;
        RECT 88.030 11.880 88.330 23.655 ;
        RECT 88.665 19.415 88.965 24.490 ;
        RECT 89.280 22.560 89.610 23.310 ;
        RECT 90.110 23.210 90.440 23.960 ;
        RECT 90.765 23.090 91.065 37.310 ;
        RECT 91.440 37.155 91.740 37.795 ;
        RECT 92.065 37.660 92.365 38.075 ;
        RECT 92.720 37.660 93.020 41.675 ;
        RECT 93.965 41.670 94.295 42.020 ;
        RECT 94.605 41.830 94.935 42.590 ;
        RECT 95.440 42.315 95.770 43.065 ;
        RECT 92.050 37.310 93.020 37.660 ;
        RECT 91.425 36.805 91.755 37.155 ;
        RECT 91.440 35.125 91.740 36.805 ;
        RECT 91.425 34.775 91.755 35.125 ;
        RECT 91.440 30.835 91.740 34.775 ;
        RECT 92.050 34.135 92.380 34.485 ;
        RECT 91.425 30.485 91.755 30.835 ;
        RECT 92.065 30.125 92.365 34.135 ;
        RECT 91.420 29.775 91.750 30.125 ;
        RECT 92.050 29.775 92.380 30.125 ;
        RECT 90.750 22.740 91.080 23.090 ;
        RECT 91.435 22.590 91.735 29.775 ;
        RECT 92.065 26.950 92.365 29.775 ;
        RECT 92.050 26.600 92.380 26.950 ;
        RECT 92.720 23.955 93.020 37.310 ;
        RECT 93.335 34.135 93.665 34.485 ;
        RECT 93.350 27.365 93.650 34.135 ;
        RECT 93.350 26.950 93.665 27.365 ;
        RECT 93.350 26.600 93.680 26.950 ;
        RECT 93.350 24.790 93.650 26.600 ;
        RECT 93.980 26.365 94.280 41.670 ;
        RECT 94.610 40.385 94.940 41.135 ;
        RECT 95.440 41.015 95.770 41.765 ;
        RECT 94.605 37.630 94.935 38.380 ;
        RECT 95.445 38.280 95.775 39.030 ;
        RECT 96.100 37.660 96.400 52.960 ;
        RECT 96.770 52.730 97.085 53.145 ;
        RECT 96.770 52.380 97.100 52.730 ;
        RECT 98.015 52.380 98.345 52.730 ;
        RECT 96.770 45.195 97.070 52.380 ;
        RECT 98.030 49.560 98.330 52.380 ;
        RECT 97.385 49.205 97.715 49.555 ;
        RECT 98.015 49.210 98.345 49.560 ;
        RECT 98.685 49.555 98.985 56.740 ;
        RECT 99.300 56.235 99.630 56.585 ;
        RECT 97.400 45.195 97.700 49.205 ;
        RECT 98.030 45.195 98.330 49.210 ;
        RECT 98.670 49.205 99.000 49.555 ;
        RECT 96.755 44.845 97.085 45.195 ;
        RECT 97.385 44.845 97.715 45.195 ;
        RECT 98.015 44.845 98.345 45.195 ;
        RECT 97.400 42.020 97.700 44.845 ;
        RECT 97.385 41.670 97.715 42.020 ;
        RECT 98.040 41.675 98.370 42.025 ;
        RECT 99.315 42.020 99.615 56.235 ;
        RECT 99.945 55.455 100.275 56.205 ;
        RECT 100.765 56.085 101.095 56.835 ;
        RECT 99.940 52.700 100.270 53.450 ;
        RECT 100.770 53.350 101.100 54.100 ;
        RECT 101.410 52.960 101.740 53.310 ;
        RECT 102.095 53.145 102.395 59.915 ;
        RECT 102.725 57.090 103.025 59.915 ;
        RECT 104.010 57.505 104.310 64.275 ;
        RECT 105.270 62.990 105.600 63.740 ;
        RECT 106.100 63.620 106.430 64.370 ;
        RECT 108.045 64.275 108.375 64.625 ;
        RECT 108.675 64.280 109.005 64.630 ;
        RECT 105.265 60.235 105.595 60.985 ;
        RECT 106.105 60.885 106.435 61.635 ;
        RECT 108.060 60.265 108.360 64.275 ;
        RECT 108.690 60.265 108.990 64.280 ;
        RECT 109.330 64.275 109.660 64.625 ;
        RECT 110.600 64.435 110.930 65.195 ;
        RECT 111.425 64.920 111.755 65.670 ;
        RECT 114.015 64.630 114.315 67.450 ;
        RECT 115.925 66.485 116.255 67.235 ;
        RECT 117.940 66.300 118.240 67.450 ;
        RECT 117.930 65.920 118.250 66.300 ;
        RECT 105.265 58.950 105.595 59.700 ;
        RECT 106.100 59.350 106.430 60.105 ;
        RECT 107.415 59.915 107.745 60.265 ;
        RECT 108.045 59.915 108.375 60.265 ;
        RECT 108.675 59.915 109.005 60.265 ;
        RECT 104.010 57.090 104.325 57.505 ;
        RECT 102.710 56.740 103.040 57.090 ;
        RECT 104.010 56.740 104.340 57.090 ;
        RECT 105.265 56.900 105.595 57.660 ;
        RECT 106.100 57.385 106.430 58.135 ;
        RECT 99.940 51.415 100.270 52.165 ;
        RECT 100.765 51.815 101.095 52.570 ;
        RECT 99.940 49.365 100.270 50.125 ;
        RECT 100.765 49.850 101.095 50.600 ;
        RECT 99.945 47.920 100.275 48.670 ;
        RECT 100.765 48.550 101.095 49.300 ;
        RECT 99.940 45.165 100.270 45.915 ;
        RECT 100.770 45.815 101.100 46.565 ;
        RECT 99.940 43.880 100.270 44.630 ;
        RECT 100.765 44.280 101.095 45.035 ;
        RECT 94.605 36.345 94.935 37.095 ;
        RECT 95.440 36.745 95.770 37.500 ;
        RECT 96.085 37.310 96.415 37.660 ;
        RECT 94.605 34.295 94.935 35.055 ;
        RECT 95.440 34.780 95.770 35.530 ;
        RECT 94.610 32.850 94.940 33.600 ;
        RECT 95.440 33.480 95.770 34.230 ;
        RECT 94.605 30.095 94.935 30.845 ;
        RECT 95.445 30.745 95.775 31.495 ;
        RECT 94.605 28.810 94.935 29.560 ;
        RECT 95.440 29.210 95.770 29.965 ;
        RECT 94.605 26.760 94.935 27.520 ;
        RECT 95.440 27.245 95.770 27.995 ;
        RECT 93.965 26.015 94.295 26.365 ;
        RECT 94.610 25.315 94.940 26.065 ;
        RECT 95.440 25.945 95.770 26.695 ;
        RECT 93.350 24.490 94.290 24.790 ;
        RECT 92.720 23.655 93.655 23.955 ;
        RECT 89.280 21.275 89.610 22.025 ;
        RECT 90.105 21.675 90.435 22.430 ;
        RECT 91.420 22.240 91.750 22.590 ;
        RECT 92.680 22.240 93.010 22.590 ;
        RECT 88.650 19.065 88.980 19.415 ;
        RECT 89.280 19.225 89.610 19.985 ;
        RECT 90.105 19.710 90.435 20.460 ;
        RECT 89.285 17.780 89.615 18.530 ;
        RECT 90.105 18.410 90.435 19.160 ;
        RECT 89.280 15.025 89.610 15.775 ;
        RECT 90.110 15.675 90.440 16.425 ;
        RECT 91.435 15.055 91.735 22.240 ;
        RECT 92.695 19.420 92.995 22.240 ;
        RECT 92.050 19.065 92.380 19.415 ;
        RECT 92.680 19.070 93.010 19.420 ;
        RECT 92.065 15.055 92.365 19.065 ;
        RECT 92.695 15.055 92.995 19.070 ;
        RECT 89.280 13.740 89.610 14.490 ;
        RECT 90.105 14.140 90.435 14.895 ;
        RECT 91.420 14.705 91.750 15.055 ;
        RECT 92.050 14.705 92.380 15.055 ;
        RECT 92.680 14.705 93.010 15.055 ;
        RECT 87.380 9.750 87.680 11.535 ;
        RECT 88.015 11.530 88.345 11.880 ;
        RECT 89.280 11.620 89.610 12.450 ;
        RECT 90.105 12.175 90.435 12.925 ;
        RECT 92.065 11.880 92.365 14.705 ;
        RECT 88.660 11.310 89.610 11.620 ;
        RECT 88.660 10.610 88.970 11.310 ;
        RECT 88.650 10.240 88.980 10.610 ;
        RECT 89.285 10.245 89.615 10.995 ;
        RECT 90.105 10.875 90.435 11.625 ;
        RECT 92.050 11.530 92.380 11.880 ;
        RECT 92.690 11.535 93.020 11.885 ;
        RECT 93.355 11.880 93.655 23.655 ;
        RECT 93.990 19.415 94.290 24.490 ;
        RECT 94.605 22.560 94.935 23.310 ;
        RECT 95.445 23.210 95.775 23.960 ;
        RECT 96.100 23.090 96.400 37.310 ;
        RECT 96.775 37.155 97.075 37.795 ;
        RECT 97.400 37.660 97.700 38.075 ;
        RECT 98.055 37.660 98.355 41.675 ;
        RECT 99.300 41.670 99.630 42.020 ;
        RECT 99.940 41.830 100.270 42.590 ;
        RECT 100.765 42.315 101.095 43.065 ;
        RECT 97.385 37.310 98.355 37.660 ;
        RECT 96.760 36.805 97.090 37.155 ;
        RECT 96.775 35.125 97.075 36.805 ;
        RECT 96.760 34.775 97.090 35.125 ;
        RECT 96.775 30.835 97.075 34.775 ;
        RECT 97.385 34.135 97.715 34.485 ;
        RECT 96.760 30.485 97.090 30.835 ;
        RECT 97.400 30.125 97.700 34.135 ;
        RECT 96.755 29.775 97.085 30.125 ;
        RECT 97.385 29.775 97.715 30.125 ;
        RECT 96.085 22.740 96.415 23.090 ;
        RECT 96.770 22.590 97.070 29.775 ;
        RECT 97.400 26.950 97.700 29.775 ;
        RECT 97.385 26.600 97.715 26.950 ;
        RECT 98.055 23.955 98.355 37.310 ;
        RECT 98.670 34.135 99.000 34.485 ;
        RECT 98.685 27.365 98.985 34.135 ;
        RECT 98.685 26.950 99.000 27.365 ;
        RECT 98.685 26.600 99.015 26.950 ;
        RECT 98.685 24.790 98.985 26.600 ;
        RECT 99.315 26.365 99.615 41.670 ;
        RECT 99.945 40.385 100.275 41.135 ;
        RECT 100.765 41.015 101.095 41.765 ;
        RECT 99.940 37.630 100.270 38.380 ;
        RECT 100.770 38.280 101.100 39.030 ;
        RECT 101.425 37.660 101.725 52.960 ;
        RECT 102.095 52.730 102.410 53.145 ;
        RECT 102.095 52.380 102.425 52.730 ;
        RECT 103.340 52.380 103.670 52.730 ;
        RECT 102.095 45.195 102.395 52.380 ;
        RECT 103.355 49.560 103.655 52.380 ;
        RECT 102.710 49.205 103.040 49.555 ;
        RECT 103.340 49.210 103.670 49.560 ;
        RECT 104.010 49.555 104.310 56.740 ;
        RECT 104.625 56.235 104.955 56.585 ;
        RECT 102.725 45.195 103.025 49.205 ;
        RECT 103.355 45.195 103.655 49.210 ;
        RECT 103.995 49.205 104.325 49.555 ;
        RECT 102.080 44.845 102.410 45.195 ;
        RECT 102.710 44.845 103.040 45.195 ;
        RECT 103.340 44.845 103.670 45.195 ;
        RECT 102.725 42.020 103.025 44.845 ;
        RECT 102.710 41.670 103.040 42.020 ;
        RECT 103.365 41.675 103.695 42.025 ;
        RECT 104.640 42.020 104.940 56.235 ;
        RECT 105.270 55.455 105.600 56.205 ;
        RECT 106.100 56.085 106.430 56.835 ;
        RECT 105.265 52.700 105.595 53.450 ;
        RECT 106.105 53.350 106.435 54.100 ;
        RECT 106.745 52.960 107.075 53.310 ;
        RECT 107.430 53.145 107.730 59.915 ;
        RECT 108.060 57.090 108.360 59.915 ;
        RECT 109.345 57.505 109.645 64.275 ;
        RECT 110.605 62.990 110.935 63.740 ;
        RECT 111.425 63.620 111.755 64.370 ;
        RECT 113.370 64.275 113.700 64.625 ;
        RECT 114.000 64.280 114.330 64.630 ;
        RECT 110.600 60.235 110.930 60.985 ;
        RECT 111.430 60.885 111.760 61.635 ;
        RECT 113.385 60.265 113.685 64.275 ;
        RECT 114.015 60.265 114.315 64.280 ;
        RECT 114.655 64.275 114.985 64.625 ;
        RECT 115.925 64.435 116.255 65.195 ;
        RECT 116.760 64.920 117.090 65.670 ;
        RECT 119.350 64.630 119.650 67.450 ;
        RECT 121.260 66.485 121.590 67.235 ;
        RECT 110.600 58.950 110.930 59.700 ;
        RECT 111.425 59.350 111.755 60.105 ;
        RECT 112.740 59.915 113.070 60.265 ;
        RECT 113.370 59.915 113.700 60.265 ;
        RECT 114.000 59.915 114.330 60.265 ;
        RECT 109.345 57.090 109.660 57.505 ;
        RECT 108.045 56.740 108.375 57.090 ;
        RECT 109.345 56.740 109.675 57.090 ;
        RECT 110.600 56.900 110.930 57.660 ;
        RECT 111.425 57.385 111.755 58.135 ;
        RECT 105.265 51.415 105.595 52.165 ;
        RECT 106.100 51.815 106.430 52.570 ;
        RECT 105.265 49.365 105.595 50.125 ;
        RECT 106.100 49.850 106.430 50.600 ;
        RECT 105.270 47.920 105.600 48.670 ;
        RECT 106.100 48.550 106.430 49.300 ;
        RECT 105.265 45.165 105.595 45.915 ;
        RECT 106.105 45.815 106.435 46.565 ;
        RECT 105.265 43.880 105.595 44.630 ;
        RECT 106.100 44.280 106.430 45.035 ;
        RECT 99.940 36.345 100.270 37.095 ;
        RECT 100.765 36.745 101.095 37.500 ;
        RECT 101.410 37.310 101.740 37.660 ;
        RECT 99.940 34.295 100.270 35.055 ;
        RECT 100.765 34.780 101.095 35.530 ;
        RECT 99.945 32.850 100.275 33.600 ;
        RECT 100.765 33.480 101.095 34.230 ;
        RECT 99.940 30.095 100.270 30.845 ;
        RECT 100.770 30.745 101.100 31.495 ;
        RECT 99.940 28.810 100.270 29.560 ;
        RECT 100.765 29.210 101.095 29.965 ;
        RECT 99.940 26.760 100.270 27.520 ;
        RECT 100.765 27.245 101.095 27.995 ;
        RECT 99.300 26.015 99.630 26.365 ;
        RECT 99.945 25.315 100.275 26.065 ;
        RECT 100.765 25.945 101.095 26.695 ;
        RECT 98.685 24.490 99.625 24.790 ;
        RECT 98.055 23.655 98.990 23.955 ;
        RECT 94.605 21.275 94.935 22.025 ;
        RECT 95.440 21.675 95.770 22.430 ;
        RECT 96.755 22.240 97.085 22.590 ;
        RECT 98.015 22.240 98.345 22.590 ;
        RECT 93.975 19.065 94.305 19.415 ;
        RECT 94.605 19.225 94.935 19.985 ;
        RECT 95.440 19.710 95.770 20.460 ;
        RECT 94.610 17.780 94.940 18.530 ;
        RECT 95.440 18.410 95.770 19.160 ;
        RECT 94.605 15.025 94.935 15.775 ;
        RECT 95.445 15.675 95.775 16.425 ;
        RECT 96.770 15.055 97.070 22.240 ;
        RECT 98.030 19.420 98.330 22.240 ;
        RECT 97.385 19.065 97.715 19.415 ;
        RECT 98.015 19.070 98.345 19.420 ;
        RECT 97.400 15.055 97.700 19.065 ;
        RECT 98.030 15.055 98.330 19.070 ;
        RECT 94.605 13.740 94.935 14.490 ;
        RECT 95.440 14.140 95.770 14.895 ;
        RECT 96.755 14.705 97.085 15.055 ;
        RECT 97.385 14.705 97.715 15.055 ;
        RECT 98.015 14.705 98.345 15.055 ;
        RECT 82.035 9.210 82.355 9.590 ;
        RECT 87.370 9.370 87.690 9.750 ;
        RECT 92.705 9.590 93.005 11.535 ;
        RECT 93.340 11.530 93.670 11.880 ;
        RECT 94.605 11.690 94.935 12.450 ;
        RECT 95.440 12.175 95.770 12.925 ;
        RECT 97.400 11.880 97.700 14.705 ;
        RECT 94.610 10.245 94.940 10.995 ;
        RECT 95.440 10.875 95.770 11.625 ;
        RECT 97.385 11.530 97.715 11.880 ;
        RECT 98.025 11.535 98.355 11.885 ;
        RECT 98.690 11.880 98.990 23.655 ;
        RECT 99.325 19.415 99.625 24.490 ;
        RECT 99.940 22.560 100.270 23.310 ;
        RECT 100.770 23.210 101.100 23.960 ;
        RECT 101.425 23.090 101.725 37.310 ;
        RECT 102.100 37.155 102.400 37.795 ;
        RECT 102.725 37.660 103.025 38.075 ;
        RECT 103.380 37.660 103.680 41.675 ;
        RECT 104.625 41.670 104.955 42.020 ;
        RECT 105.265 41.830 105.595 42.590 ;
        RECT 106.100 42.315 106.430 43.065 ;
        RECT 102.710 37.310 103.680 37.660 ;
        RECT 102.085 36.805 102.415 37.155 ;
        RECT 102.100 35.125 102.400 36.805 ;
        RECT 102.085 34.775 102.415 35.125 ;
        RECT 102.100 30.835 102.400 34.775 ;
        RECT 102.710 34.135 103.040 34.485 ;
        RECT 102.085 30.485 102.415 30.835 ;
        RECT 102.725 30.125 103.025 34.135 ;
        RECT 102.080 29.775 102.410 30.125 ;
        RECT 102.710 29.775 103.040 30.125 ;
        RECT 101.410 22.740 101.740 23.090 ;
        RECT 102.095 22.590 102.395 29.775 ;
        RECT 102.725 26.950 103.025 29.775 ;
        RECT 102.710 26.600 103.040 26.950 ;
        RECT 103.380 23.955 103.680 37.310 ;
        RECT 103.995 34.135 104.325 34.485 ;
        RECT 104.010 27.365 104.310 34.135 ;
        RECT 104.010 26.950 104.325 27.365 ;
        RECT 104.010 26.600 104.340 26.950 ;
        RECT 104.010 24.790 104.310 26.600 ;
        RECT 104.640 26.365 104.940 41.670 ;
        RECT 105.270 40.385 105.600 41.135 ;
        RECT 106.100 41.015 106.430 41.765 ;
        RECT 105.265 37.630 105.595 38.380 ;
        RECT 106.105 38.280 106.435 39.030 ;
        RECT 106.760 37.660 107.060 52.960 ;
        RECT 107.430 52.730 107.745 53.145 ;
        RECT 107.430 52.380 107.760 52.730 ;
        RECT 108.675 52.380 109.005 52.730 ;
        RECT 107.430 45.195 107.730 52.380 ;
        RECT 108.690 49.560 108.990 52.380 ;
        RECT 108.045 49.205 108.375 49.555 ;
        RECT 108.675 49.210 109.005 49.560 ;
        RECT 109.345 49.555 109.645 56.740 ;
        RECT 109.960 56.235 110.290 56.585 ;
        RECT 108.060 45.195 108.360 49.205 ;
        RECT 108.690 45.195 108.990 49.210 ;
        RECT 109.330 49.205 109.660 49.555 ;
        RECT 107.415 44.845 107.745 45.195 ;
        RECT 108.045 44.845 108.375 45.195 ;
        RECT 108.675 44.845 109.005 45.195 ;
        RECT 108.060 42.020 108.360 44.845 ;
        RECT 108.045 41.670 108.375 42.020 ;
        RECT 108.700 41.675 109.030 42.025 ;
        RECT 109.975 42.020 110.275 56.235 ;
        RECT 110.605 55.455 110.935 56.205 ;
        RECT 111.425 56.085 111.755 56.835 ;
        RECT 110.600 52.700 110.930 53.450 ;
        RECT 111.430 53.350 111.760 54.100 ;
        RECT 112.070 52.960 112.400 53.310 ;
        RECT 112.755 53.145 113.055 59.915 ;
        RECT 113.385 57.090 113.685 59.915 ;
        RECT 114.670 57.505 114.970 64.275 ;
        RECT 115.930 62.990 116.260 63.740 ;
        RECT 116.760 63.620 117.090 64.370 ;
        RECT 118.705 64.275 119.035 64.625 ;
        RECT 119.335 64.280 119.665 64.630 ;
        RECT 115.925 60.235 116.255 60.985 ;
        RECT 116.765 60.885 117.095 61.635 ;
        RECT 118.720 60.265 119.020 64.275 ;
        RECT 119.350 60.265 119.650 64.280 ;
        RECT 119.990 64.275 120.320 64.625 ;
        RECT 121.260 64.435 121.590 65.195 ;
        RECT 115.925 58.950 116.255 59.700 ;
        RECT 116.760 59.350 117.090 60.105 ;
        RECT 118.075 59.915 118.405 60.265 ;
        RECT 118.705 59.915 119.035 60.265 ;
        RECT 119.335 59.915 119.665 60.265 ;
        RECT 114.670 57.090 114.985 57.505 ;
        RECT 113.370 56.740 113.700 57.090 ;
        RECT 114.670 56.740 115.000 57.090 ;
        RECT 115.925 56.900 116.255 57.660 ;
        RECT 116.760 57.385 117.090 58.135 ;
        RECT 110.600 51.415 110.930 52.165 ;
        RECT 111.425 51.815 111.755 52.570 ;
        RECT 110.600 49.365 110.930 50.125 ;
        RECT 111.425 49.850 111.755 50.600 ;
        RECT 110.605 47.920 110.935 48.670 ;
        RECT 111.425 48.550 111.755 49.300 ;
        RECT 110.600 45.165 110.930 45.915 ;
        RECT 111.430 45.815 111.760 46.565 ;
        RECT 110.600 43.880 110.930 44.630 ;
        RECT 111.425 44.280 111.755 45.035 ;
        RECT 105.265 36.345 105.595 37.095 ;
        RECT 106.100 36.745 106.430 37.500 ;
        RECT 106.745 37.310 107.075 37.660 ;
        RECT 105.265 34.295 105.595 35.055 ;
        RECT 106.100 34.780 106.430 35.530 ;
        RECT 105.270 32.850 105.600 33.600 ;
        RECT 106.100 33.480 106.430 34.230 ;
        RECT 105.265 30.095 105.595 30.845 ;
        RECT 106.105 30.745 106.435 31.495 ;
        RECT 105.265 28.810 105.595 29.560 ;
        RECT 106.100 29.210 106.430 29.965 ;
        RECT 105.265 26.760 105.595 27.520 ;
        RECT 106.100 27.245 106.430 27.995 ;
        RECT 104.625 26.015 104.955 26.365 ;
        RECT 105.270 25.315 105.600 26.065 ;
        RECT 106.100 25.945 106.430 26.695 ;
        RECT 104.010 24.490 104.950 24.790 ;
        RECT 103.380 23.655 104.315 23.955 ;
        RECT 99.940 21.275 100.270 22.025 ;
        RECT 100.765 21.675 101.095 22.430 ;
        RECT 102.080 22.240 102.410 22.590 ;
        RECT 103.340 22.240 103.670 22.590 ;
        RECT 99.310 19.065 99.640 19.415 ;
        RECT 99.940 19.225 100.270 19.985 ;
        RECT 100.765 19.710 101.095 20.460 ;
        RECT 99.945 17.780 100.275 18.530 ;
        RECT 100.765 18.410 101.095 19.160 ;
        RECT 99.940 15.025 100.270 15.775 ;
        RECT 100.770 15.675 101.100 16.425 ;
        RECT 102.095 15.055 102.395 22.240 ;
        RECT 103.355 19.420 103.655 22.240 ;
        RECT 102.710 19.065 103.040 19.415 ;
        RECT 103.340 19.070 103.670 19.420 ;
        RECT 102.725 15.055 103.025 19.065 ;
        RECT 103.355 15.055 103.655 19.070 ;
        RECT 99.940 13.740 100.270 14.490 ;
        RECT 100.765 14.140 101.095 14.895 ;
        RECT 102.080 14.705 102.410 15.055 ;
        RECT 102.710 14.705 103.040 15.055 ;
        RECT 103.340 14.705 103.670 15.055 ;
        RECT 98.040 9.750 98.340 11.535 ;
        RECT 98.675 11.530 99.005 11.880 ;
        RECT 99.940 11.620 100.270 12.450 ;
        RECT 100.765 12.175 101.095 12.925 ;
        RECT 102.725 11.880 103.025 14.705 ;
        RECT 99.320 11.310 100.270 11.620 ;
        RECT 99.320 10.610 99.630 11.310 ;
        RECT 99.310 10.240 99.640 10.610 ;
        RECT 99.945 10.245 100.275 10.995 ;
        RECT 100.765 10.875 101.095 11.625 ;
        RECT 102.710 11.530 103.040 11.880 ;
        RECT 103.350 11.535 103.680 11.885 ;
        RECT 104.015 11.880 104.315 23.655 ;
        RECT 104.650 19.415 104.950 24.490 ;
        RECT 105.265 22.560 105.595 23.310 ;
        RECT 106.105 23.210 106.435 23.960 ;
        RECT 106.760 23.090 107.060 37.310 ;
        RECT 107.435 37.155 107.735 37.795 ;
        RECT 108.060 37.660 108.360 38.075 ;
        RECT 108.715 37.660 109.015 41.675 ;
        RECT 109.960 41.670 110.290 42.020 ;
        RECT 110.600 41.830 110.930 42.590 ;
        RECT 111.425 42.315 111.755 43.065 ;
        RECT 108.045 37.310 109.015 37.660 ;
        RECT 107.420 36.805 107.750 37.155 ;
        RECT 107.435 35.125 107.735 36.805 ;
        RECT 107.420 34.775 107.750 35.125 ;
        RECT 107.435 30.835 107.735 34.775 ;
        RECT 108.045 34.135 108.375 34.485 ;
        RECT 107.420 30.485 107.750 30.835 ;
        RECT 108.060 30.125 108.360 34.135 ;
        RECT 107.415 29.775 107.745 30.125 ;
        RECT 108.045 29.775 108.375 30.125 ;
        RECT 106.745 22.740 107.075 23.090 ;
        RECT 107.430 22.590 107.730 29.775 ;
        RECT 108.060 26.950 108.360 29.775 ;
        RECT 108.045 26.600 108.375 26.950 ;
        RECT 108.715 23.955 109.015 37.310 ;
        RECT 109.330 34.135 109.660 34.485 ;
        RECT 109.345 27.365 109.645 34.135 ;
        RECT 109.345 26.950 109.660 27.365 ;
        RECT 109.345 26.600 109.675 26.950 ;
        RECT 109.345 24.790 109.645 26.600 ;
        RECT 109.975 26.365 110.275 41.670 ;
        RECT 110.605 40.385 110.935 41.135 ;
        RECT 111.425 41.015 111.755 41.765 ;
        RECT 110.600 37.630 110.930 38.380 ;
        RECT 111.430 38.280 111.760 39.030 ;
        RECT 112.085 37.660 112.385 52.960 ;
        RECT 112.755 52.730 113.070 53.145 ;
        RECT 112.755 52.380 113.085 52.730 ;
        RECT 114.000 52.380 114.330 52.730 ;
        RECT 112.755 45.195 113.055 52.380 ;
        RECT 114.015 49.560 114.315 52.380 ;
        RECT 113.370 49.205 113.700 49.555 ;
        RECT 114.000 49.210 114.330 49.560 ;
        RECT 114.670 49.555 114.970 56.740 ;
        RECT 115.285 56.235 115.615 56.585 ;
        RECT 113.385 45.195 113.685 49.205 ;
        RECT 114.015 45.195 114.315 49.210 ;
        RECT 114.655 49.205 114.985 49.555 ;
        RECT 112.740 44.845 113.070 45.195 ;
        RECT 113.370 44.845 113.700 45.195 ;
        RECT 114.000 44.845 114.330 45.195 ;
        RECT 113.385 42.020 113.685 44.845 ;
        RECT 113.370 41.670 113.700 42.020 ;
        RECT 114.025 41.675 114.355 42.025 ;
        RECT 115.300 42.020 115.600 56.235 ;
        RECT 115.930 55.455 116.260 56.205 ;
        RECT 116.760 56.085 117.090 56.835 ;
        RECT 115.925 52.700 116.255 53.450 ;
        RECT 116.765 53.350 117.095 54.100 ;
        RECT 117.405 52.960 117.735 53.310 ;
        RECT 118.090 53.145 118.390 59.915 ;
        RECT 118.720 57.090 119.020 59.915 ;
        RECT 120.005 57.505 120.305 64.275 ;
        RECT 121.265 62.990 121.595 63.740 ;
        RECT 121.260 60.235 121.590 60.985 ;
        RECT 121.260 58.950 121.590 59.700 ;
        RECT 120.005 57.090 120.320 57.505 ;
        RECT 118.705 56.740 119.035 57.090 ;
        RECT 120.005 56.740 120.335 57.090 ;
        RECT 121.260 56.900 121.590 57.660 ;
        RECT 115.925 51.415 116.255 52.165 ;
        RECT 116.760 51.815 117.090 52.570 ;
        RECT 115.925 49.365 116.255 50.125 ;
        RECT 116.760 49.850 117.090 50.600 ;
        RECT 115.930 47.920 116.260 48.670 ;
        RECT 116.760 48.550 117.090 49.300 ;
        RECT 115.925 45.165 116.255 45.915 ;
        RECT 116.765 45.815 117.095 46.565 ;
        RECT 115.925 43.880 116.255 44.630 ;
        RECT 116.760 44.280 117.090 45.035 ;
        RECT 110.600 36.345 110.930 37.095 ;
        RECT 111.425 36.745 111.755 37.500 ;
        RECT 112.070 37.310 112.400 37.660 ;
        RECT 110.600 34.295 110.930 35.055 ;
        RECT 111.425 34.780 111.755 35.530 ;
        RECT 110.605 32.850 110.935 33.600 ;
        RECT 111.425 33.480 111.755 34.230 ;
        RECT 110.600 30.095 110.930 30.845 ;
        RECT 111.430 30.745 111.760 31.495 ;
        RECT 110.600 28.810 110.930 29.560 ;
        RECT 111.425 29.210 111.755 29.965 ;
        RECT 110.600 26.760 110.930 27.520 ;
        RECT 111.425 27.245 111.755 27.995 ;
        RECT 109.960 26.015 110.290 26.365 ;
        RECT 110.605 25.315 110.935 26.065 ;
        RECT 111.425 25.945 111.755 26.695 ;
        RECT 109.345 24.490 110.285 24.790 ;
        RECT 108.715 23.655 109.650 23.955 ;
        RECT 105.265 21.275 105.595 22.025 ;
        RECT 106.100 21.675 106.430 22.430 ;
        RECT 107.415 22.240 107.745 22.590 ;
        RECT 108.675 22.240 109.005 22.590 ;
        RECT 104.635 19.065 104.965 19.415 ;
        RECT 105.265 19.225 105.595 19.985 ;
        RECT 106.100 19.710 106.430 20.460 ;
        RECT 105.270 17.780 105.600 18.530 ;
        RECT 106.100 18.410 106.430 19.160 ;
        RECT 105.265 15.025 105.595 15.775 ;
        RECT 106.105 15.675 106.435 16.425 ;
        RECT 107.430 15.055 107.730 22.240 ;
        RECT 108.690 19.420 108.990 22.240 ;
        RECT 108.045 19.065 108.375 19.415 ;
        RECT 108.675 19.070 109.005 19.420 ;
        RECT 108.060 15.055 108.360 19.065 ;
        RECT 108.690 15.055 108.990 19.070 ;
        RECT 105.265 13.740 105.595 14.490 ;
        RECT 106.100 14.140 106.430 14.895 ;
        RECT 107.415 14.705 107.745 15.055 ;
        RECT 108.045 14.705 108.375 15.055 ;
        RECT 108.675 14.705 109.005 15.055 ;
        RECT 92.695 9.210 93.015 9.590 ;
        RECT 98.030 9.370 98.350 9.750 ;
        RECT 103.365 9.590 103.665 11.535 ;
        RECT 104.000 11.530 104.330 11.880 ;
        RECT 105.265 11.690 105.595 12.450 ;
        RECT 106.100 12.175 106.430 12.925 ;
        RECT 108.060 11.880 108.360 14.705 ;
        RECT 105.270 10.245 105.600 10.995 ;
        RECT 106.100 10.875 106.430 11.625 ;
        RECT 108.045 11.530 108.375 11.880 ;
        RECT 108.685 11.535 109.015 11.885 ;
        RECT 109.350 11.880 109.650 23.655 ;
        RECT 109.985 19.415 110.285 24.490 ;
        RECT 110.600 22.560 110.930 23.310 ;
        RECT 111.430 23.210 111.760 23.960 ;
        RECT 112.085 23.090 112.385 37.310 ;
        RECT 112.760 37.155 113.060 37.795 ;
        RECT 113.385 37.660 113.685 38.075 ;
        RECT 114.040 37.660 114.340 41.675 ;
        RECT 115.285 41.670 115.615 42.020 ;
        RECT 115.925 41.830 116.255 42.590 ;
        RECT 116.760 42.315 117.090 43.065 ;
        RECT 113.370 37.310 114.340 37.660 ;
        RECT 112.745 36.805 113.075 37.155 ;
        RECT 112.760 35.125 113.060 36.805 ;
        RECT 112.745 34.775 113.075 35.125 ;
        RECT 112.760 30.835 113.060 34.775 ;
        RECT 113.370 34.135 113.700 34.485 ;
        RECT 112.745 30.485 113.075 30.835 ;
        RECT 113.385 30.125 113.685 34.135 ;
        RECT 112.740 29.775 113.070 30.125 ;
        RECT 113.370 29.775 113.700 30.125 ;
        RECT 112.070 22.740 112.400 23.090 ;
        RECT 112.755 22.590 113.055 29.775 ;
        RECT 113.385 26.950 113.685 29.775 ;
        RECT 113.370 26.600 113.700 26.950 ;
        RECT 114.040 23.955 114.340 37.310 ;
        RECT 114.655 34.135 114.985 34.485 ;
        RECT 114.670 27.365 114.970 34.135 ;
        RECT 114.670 26.950 114.985 27.365 ;
        RECT 114.670 26.600 115.000 26.950 ;
        RECT 114.670 24.790 114.970 26.600 ;
        RECT 115.300 26.365 115.600 41.670 ;
        RECT 115.930 40.385 116.260 41.135 ;
        RECT 116.760 41.015 117.090 41.765 ;
        RECT 115.925 37.630 116.255 38.380 ;
        RECT 116.765 38.280 117.095 39.030 ;
        RECT 117.420 37.660 117.720 52.960 ;
        RECT 118.090 52.730 118.405 53.145 ;
        RECT 118.090 52.380 118.420 52.730 ;
        RECT 119.335 52.380 119.665 52.730 ;
        RECT 118.090 45.195 118.390 52.380 ;
        RECT 119.350 49.560 119.650 52.380 ;
        RECT 118.705 49.205 119.035 49.555 ;
        RECT 119.335 49.210 119.665 49.560 ;
        RECT 120.005 49.555 120.305 56.740 ;
        RECT 120.620 56.235 120.950 56.585 ;
        RECT 118.720 45.195 119.020 49.205 ;
        RECT 119.350 45.195 119.650 49.210 ;
        RECT 119.990 49.205 120.320 49.555 ;
        RECT 118.075 44.845 118.405 45.195 ;
        RECT 118.705 44.845 119.035 45.195 ;
        RECT 119.335 44.845 119.665 45.195 ;
        RECT 118.720 42.020 119.020 44.845 ;
        RECT 118.705 41.670 119.035 42.020 ;
        RECT 119.360 41.675 119.690 42.025 ;
        RECT 120.635 42.020 120.935 56.235 ;
        RECT 121.265 55.455 121.595 56.205 ;
        RECT 121.260 52.700 121.590 53.450 ;
        RECT 121.260 51.415 121.590 52.165 ;
        RECT 121.260 49.365 121.590 50.125 ;
        RECT 121.265 47.920 121.595 48.670 ;
        RECT 121.260 45.165 121.590 45.915 ;
        RECT 121.260 43.880 121.590 44.630 ;
        RECT 115.925 36.345 116.255 37.095 ;
        RECT 116.760 36.745 117.090 37.500 ;
        RECT 117.405 37.310 117.735 37.660 ;
        RECT 115.925 34.295 116.255 35.055 ;
        RECT 116.760 34.780 117.090 35.530 ;
        RECT 115.930 32.850 116.260 33.600 ;
        RECT 116.760 33.480 117.090 34.230 ;
        RECT 115.925 30.095 116.255 30.845 ;
        RECT 116.765 30.745 117.095 31.495 ;
        RECT 115.925 28.810 116.255 29.560 ;
        RECT 116.760 29.210 117.090 29.965 ;
        RECT 115.925 26.760 116.255 27.520 ;
        RECT 116.760 27.245 117.090 27.995 ;
        RECT 115.285 26.015 115.615 26.365 ;
        RECT 115.930 25.315 116.260 26.065 ;
        RECT 116.760 25.945 117.090 26.695 ;
        RECT 114.670 24.490 115.610 24.790 ;
        RECT 114.040 23.655 114.975 23.955 ;
        RECT 110.600 21.275 110.930 22.025 ;
        RECT 111.425 21.675 111.755 22.430 ;
        RECT 112.740 22.240 113.070 22.590 ;
        RECT 114.000 22.240 114.330 22.590 ;
        RECT 109.970 19.065 110.300 19.415 ;
        RECT 110.600 19.225 110.930 19.985 ;
        RECT 111.425 19.710 111.755 20.460 ;
        RECT 110.605 17.780 110.935 18.530 ;
        RECT 111.425 18.410 111.755 19.160 ;
        RECT 110.600 15.025 110.930 15.775 ;
        RECT 111.430 15.675 111.760 16.425 ;
        RECT 112.755 15.055 113.055 22.240 ;
        RECT 114.015 19.420 114.315 22.240 ;
        RECT 113.370 19.065 113.700 19.415 ;
        RECT 114.000 19.070 114.330 19.420 ;
        RECT 113.385 15.055 113.685 19.065 ;
        RECT 114.015 15.055 114.315 19.070 ;
        RECT 110.600 13.740 110.930 14.490 ;
        RECT 111.425 14.140 111.755 14.895 ;
        RECT 112.740 14.705 113.070 15.055 ;
        RECT 113.370 14.705 113.700 15.055 ;
        RECT 114.000 14.705 114.330 15.055 ;
        RECT 108.700 9.750 109.000 11.535 ;
        RECT 109.335 11.530 109.665 11.880 ;
        RECT 110.600 11.620 110.930 12.450 ;
        RECT 111.425 12.175 111.755 12.925 ;
        RECT 113.385 11.880 113.685 14.705 ;
        RECT 109.980 11.310 110.930 11.620 ;
        RECT 109.980 10.610 110.290 11.310 ;
        RECT 109.970 10.240 110.300 10.610 ;
        RECT 110.605 10.245 110.935 10.995 ;
        RECT 111.425 10.875 111.755 11.625 ;
        RECT 113.370 11.530 113.700 11.880 ;
        RECT 114.010 11.535 114.340 11.885 ;
        RECT 114.675 11.880 114.975 23.655 ;
        RECT 115.310 19.415 115.610 24.490 ;
        RECT 115.925 22.560 116.255 23.310 ;
        RECT 116.765 23.210 117.095 23.960 ;
        RECT 117.420 23.090 117.720 37.310 ;
        RECT 118.095 37.155 118.395 37.795 ;
        RECT 118.720 37.660 119.020 38.075 ;
        RECT 119.375 37.660 119.675 41.675 ;
        RECT 120.620 41.670 120.950 42.020 ;
        RECT 121.260 41.830 121.590 42.590 ;
        RECT 118.705 37.310 119.675 37.660 ;
        RECT 118.080 36.805 118.410 37.155 ;
        RECT 118.095 35.125 118.395 36.805 ;
        RECT 118.080 34.775 118.410 35.125 ;
        RECT 118.095 30.835 118.395 34.775 ;
        RECT 118.705 34.135 119.035 34.485 ;
        RECT 118.080 30.485 118.410 30.835 ;
        RECT 118.720 30.125 119.020 34.135 ;
        RECT 118.075 29.775 118.405 30.125 ;
        RECT 118.705 29.775 119.035 30.125 ;
        RECT 117.405 22.740 117.735 23.090 ;
        RECT 118.090 22.590 118.390 29.775 ;
        RECT 118.720 26.950 119.020 29.775 ;
        RECT 118.705 26.600 119.035 26.950 ;
        RECT 119.375 23.955 119.675 37.310 ;
        RECT 119.990 34.135 120.320 34.485 ;
        RECT 120.005 27.365 120.305 34.135 ;
        RECT 120.005 26.950 120.320 27.365 ;
        RECT 120.005 26.600 120.335 26.950 ;
        RECT 120.005 24.790 120.305 26.600 ;
        RECT 120.635 26.365 120.935 41.670 ;
        RECT 121.265 40.385 121.595 41.135 ;
        RECT 121.260 37.630 121.590 38.380 ;
        RECT 121.260 36.345 121.590 37.095 ;
        RECT 121.260 34.295 121.590 35.055 ;
        RECT 121.265 32.850 121.595 33.600 ;
        RECT 121.260 30.095 121.590 30.845 ;
        RECT 121.260 28.810 121.590 29.560 ;
        RECT 121.260 26.760 121.590 27.520 ;
        RECT 120.620 26.015 120.950 26.365 ;
        RECT 121.265 25.315 121.595 26.065 ;
        RECT 120.005 24.490 120.945 24.790 ;
        RECT 119.375 23.655 120.310 23.955 ;
        RECT 115.925 21.275 116.255 22.025 ;
        RECT 116.760 21.675 117.090 22.430 ;
        RECT 118.075 22.240 118.405 22.590 ;
        RECT 119.335 22.240 119.665 22.590 ;
        RECT 115.295 19.065 115.625 19.415 ;
        RECT 115.925 19.225 116.255 19.985 ;
        RECT 116.760 19.710 117.090 20.460 ;
        RECT 115.930 17.780 116.260 18.530 ;
        RECT 116.760 18.410 117.090 19.160 ;
        RECT 115.925 15.025 116.255 15.775 ;
        RECT 116.765 15.675 117.095 16.425 ;
        RECT 118.090 15.055 118.390 22.240 ;
        RECT 119.350 19.420 119.650 22.240 ;
        RECT 118.705 19.065 119.035 19.415 ;
        RECT 119.335 19.070 119.665 19.420 ;
        RECT 118.720 15.055 119.020 19.065 ;
        RECT 119.350 15.055 119.650 19.070 ;
        RECT 115.925 13.740 116.255 14.490 ;
        RECT 116.760 14.140 117.090 14.895 ;
        RECT 118.075 14.705 118.405 15.055 ;
        RECT 118.705 14.705 119.035 15.055 ;
        RECT 119.335 14.705 119.665 15.055 ;
        RECT 103.355 9.210 103.675 9.590 ;
        RECT 108.690 9.370 109.010 9.750 ;
        RECT 114.025 9.590 114.325 11.535 ;
        RECT 114.660 11.530 114.990 11.880 ;
        RECT 115.925 11.690 116.255 12.450 ;
        RECT 116.760 12.175 117.090 12.925 ;
        RECT 118.720 11.880 119.020 14.705 ;
        RECT 115.930 10.245 116.260 10.995 ;
        RECT 116.760 10.875 117.090 11.625 ;
        RECT 118.705 11.530 119.035 11.880 ;
        RECT 119.345 11.535 119.675 11.885 ;
        RECT 120.010 11.880 120.310 23.655 ;
        RECT 120.645 19.415 120.945 24.490 ;
        RECT 121.260 22.560 121.590 23.310 ;
        RECT 121.260 21.275 121.590 22.025 ;
        RECT 120.630 19.065 120.960 19.415 ;
        RECT 121.260 19.225 121.590 19.985 ;
        RECT 121.265 17.780 121.595 18.530 ;
        RECT 121.260 15.025 121.590 15.775 ;
        RECT 121.260 13.740 121.590 14.490 ;
        RECT 119.360 9.750 119.660 11.535 ;
        RECT 119.995 11.530 120.325 11.880 ;
        RECT 121.260 11.620 121.590 12.450 ;
        RECT 120.640 11.310 121.590 11.620 ;
        RECT 120.640 10.610 120.950 11.310 ;
        RECT 120.630 10.240 120.960 10.610 ;
        RECT 121.265 10.245 121.595 10.995 ;
        RECT 114.015 9.210 114.335 9.590 ;
        RECT 119.350 9.370 119.670 9.750 ;
      LAYER met4 ;
        RECT 44.080 73.725 44.410 73.740 ;
        RECT 54.740 73.725 55.070 73.740 ;
        RECT 65.400 73.725 65.730 73.740 ;
        RECT 44.080 73.425 65.730 73.725 ;
        RECT 44.080 73.410 44.410 73.425 ;
        RECT 54.740 73.410 55.070 73.425 ;
        RECT 65.400 73.410 65.730 73.425 ;
        RECT 86.720 73.725 87.050 73.740 ;
        RECT 97.380 73.725 97.710 73.740 ;
        RECT 108.040 73.725 108.370 73.740 ;
        RECT 86.720 73.425 108.370 73.725 ;
        RECT 86.720 73.410 87.050 73.425 ;
        RECT 97.380 73.410 97.710 73.425 ;
        RECT 108.040 73.410 108.370 73.425 ;
        RECT 38.625 69.250 39.805 70.430 ;
        RECT 49.285 69.250 50.465 70.430 ;
        RECT 59.945 69.250 61.125 70.430 ;
        RECT 70.605 69.250 71.785 70.430 ;
        RECT 81.265 69.250 82.445 70.430 ;
        RECT 91.925 69.250 93.105 70.430 ;
        RECT 102.585 69.250 103.765 70.430 ;
        RECT 113.245 69.250 114.425 70.430 ;
        RECT 29.735 68.825 30.935 68.840 ;
        RECT 31.485 68.825 31.815 68.840 ;
        RECT 36.805 68.825 37.135 68.840 ;
        RECT 48.095 68.825 48.425 68.840 ;
        RECT 58.125 68.825 58.455 68.840 ;
        RECT 69.415 68.825 69.745 68.840 ;
        RECT 79.445 68.825 79.775 68.840 ;
        RECT 90.735 68.825 91.065 68.840 ;
        RECT 100.765 68.825 101.095 68.840 ;
        RECT 112.055 68.825 112.385 68.840 ;
        RECT 122.090 68.825 122.420 68.840 ;
        RECT 29.705 68.525 127.180 68.825 ;
        RECT 29.735 68.510 30.935 68.525 ;
        RECT 31.485 68.510 31.815 68.525 ;
        RECT 36.805 68.510 37.135 68.525 ;
        RECT 48.095 68.510 48.425 68.525 ;
        RECT 58.125 68.510 58.455 68.525 ;
        RECT 69.415 68.510 69.745 68.525 ;
        RECT 79.445 68.510 79.775 68.525 ;
        RECT 90.735 68.510 91.065 68.525 ;
        RECT 100.765 68.510 101.095 68.525 ;
        RECT 112.055 68.510 112.385 68.525 ;
        RECT 122.090 68.510 122.420 68.525 ;
        RECT 29.735 68.180 30.935 68.195 ;
        RECT 35.980 68.180 36.310 68.195 ;
        RECT 41.305 68.180 41.635 68.195 ;
        RECT 46.640 68.180 46.970 68.195 ;
        RECT 51.965 68.180 52.295 68.195 ;
        RECT 57.300 68.180 57.630 68.195 ;
        RECT 62.625 68.180 62.955 68.195 ;
        RECT 67.960 68.180 68.290 68.195 ;
        RECT 73.285 68.180 73.615 68.195 ;
        RECT 78.620 68.180 78.950 68.195 ;
        RECT 83.945 68.180 84.275 68.195 ;
        RECT 89.280 68.180 89.610 68.195 ;
        RECT 94.605 68.180 94.935 68.195 ;
        RECT 99.940 68.180 100.270 68.195 ;
        RECT 105.265 68.180 105.595 68.195 ;
        RECT 110.600 68.180 110.930 68.195 ;
        RECT 115.925 68.180 116.255 68.195 ;
        RECT 121.260 68.180 121.590 68.195 ;
        RECT 126.585 68.180 126.915 68.195 ;
        RECT 29.705 67.880 127.180 68.180 ;
        RECT 29.735 67.865 30.935 67.880 ;
        RECT 35.980 67.865 36.310 67.880 ;
        RECT 41.305 67.865 41.635 67.880 ;
        RECT 46.640 67.865 46.970 67.880 ;
        RECT 51.965 67.865 52.295 67.880 ;
        RECT 57.300 67.865 57.630 67.880 ;
        RECT 62.625 67.865 62.955 67.880 ;
        RECT 67.960 67.865 68.290 67.880 ;
        RECT 73.285 67.865 73.615 67.880 ;
        RECT 78.620 67.865 78.950 67.880 ;
        RECT 83.945 67.865 84.275 67.880 ;
        RECT 89.280 67.865 89.610 67.880 ;
        RECT 94.605 67.865 94.935 67.880 ;
        RECT 99.940 67.865 100.270 67.880 ;
        RECT 105.265 67.865 105.595 67.880 ;
        RECT 110.600 67.865 110.930 67.880 ;
        RECT 115.925 67.865 116.255 67.880 ;
        RECT 121.260 67.865 121.590 67.880 ;
        RECT 126.585 67.865 126.915 67.880 ;
        RECT 29.735 67.535 30.935 67.550 ;
        RECT 31.480 67.535 31.810 67.550 ;
        RECT 36.805 67.535 37.135 67.550 ;
        RECT 45.775 67.535 46.105 67.550 ;
        RECT 58.125 67.535 58.455 67.550 ;
        RECT 67.095 67.535 67.425 67.550 ;
        RECT 79.445 67.535 79.775 67.550 ;
        RECT 88.415 67.535 88.745 67.550 ;
        RECT 100.765 67.535 101.095 67.550 ;
        RECT 109.735 67.535 110.065 67.550 ;
        RECT 122.085 67.535 122.415 67.550 ;
        RECT 29.705 67.235 127.180 67.535 ;
        RECT 29.735 67.220 30.935 67.235 ;
        RECT 31.480 67.220 31.810 67.235 ;
        RECT 36.805 67.220 37.135 67.235 ;
        RECT 45.775 67.220 46.105 67.235 ;
        RECT 58.125 67.220 58.455 67.235 ;
        RECT 67.095 67.220 67.425 67.235 ;
        RECT 79.445 67.220 79.775 67.235 ;
        RECT 88.415 67.220 88.745 67.235 ;
        RECT 100.765 67.220 101.095 67.235 ;
        RECT 109.735 67.220 110.065 67.235 ;
        RECT 122.085 67.220 122.415 67.235 ;
        RECT 29.735 66.890 30.935 66.905 ;
        RECT 35.980 66.890 36.310 66.905 ;
        RECT 41.305 66.890 41.635 66.905 ;
        RECT 46.640 66.890 46.970 66.905 ;
        RECT 51.965 66.890 52.295 66.905 ;
        RECT 57.300 66.890 57.630 66.905 ;
        RECT 62.625 66.890 62.955 66.905 ;
        RECT 67.960 66.890 68.290 66.905 ;
        RECT 73.285 66.890 73.615 66.905 ;
        RECT 78.620 66.890 78.950 66.905 ;
        RECT 83.945 66.890 84.275 66.905 ;
        RECT 89.280 66.890 89.610 66.905 ;
        RECT 94.605 66.890 94.935 66.905 ;
        RECT 99.940 66.890 100.270 66.905 ;
        RECT 105.265 66.890 105.595 66.905 ;
        RECT 110.600 66.890 110.930 66.905 ;
        RECT 115.925 66.890 116.255 66.905 ;
        RECT 121.260 66.890 121.590 66.905 ;
        RECT 126.585 66.890 126.915 66.905 ;
        RECT 29.705 66.590 127.180 66.890 ;
        RECT 29.735 66.575 30.935 66.590 ;
        RECT 35.980 66.575 36.310 66.590 ;
        RECT 41.305 66.575 41.635 66.590 ;
        RECT 46.640 66.575 46.970 66.590 ;
        RECT 51.965 66.575 52.295 66.590 ;
        RECT 57.300 66.575 57.630 66.590 ;
        RECT 62.625 66.575 62.955 66.590 ;
        RECT 67.960 66.575 68.290 66.590 ;
        RECT 73.285 66.575 73.615 66.590 ;
        RECT 78.620 66.575 78.950 66.590 ;
        RECT 83.945 66.575 84.275 66.590 ;
        RECT 89.280 66.575 89.610 66.590 ;
        RECT 94.605 66.575 94.935 66.590 ;
        RECT 99.940 66.575 100.270 66.590 ;
        RECT 105.265 66.575 105.595 66.590 ;
        RECT 110.600 66.575 110.930 66.590 ;
        RECT 115.925 66.575 116.255 66.590 ;
        RECT 121.260 66.575 121.590 66.590 ;
        RECT 126.585 66.575 126.915 66.590 ;
        RECT 37.970 66.260 38.300 66.275 ;
        RECT 43.305 66.260 43.635 66.275 ;
        RECT 48.630 66.260 48.960 66.275 ;
        RECT 59.290 66.260 59.620 66.275 ;
        RECT 64.625 66.260 64.955 66.275 ;
        RECT 69.950 66.260 70.280 66.275 ;
        RECT 75.285 66.260 75.615 66.275 ;
        RECT 77.585 66.260 77.915 66.275 ;
        RECT 37.970 65.960 49.400 66.260 ;
        RECT 59.290 65.960 70.720 66.260 ;
        RECT 74.845 65.960 75.615 66.260 ;
        RECT 77.145 65.960 77.915 66.260 ;
        RECT 37.970 65.945 38.300 65.960 ;
        RECT 43.305 65.945 43.635 65.960 ;
        RECT 48.630 65.945 48.960 65.960 ;
        RECT 59.290 65.945 59.620 65.960 ;
        RECT 64.625 65.945 64.955 65.960 ;
        RECT 69.950 65.945 70.280 65.960 ;
        RECT 75.285 65.945 75.615 65.960 ;
        RECT 77.585 65.945 77.915 65.960 ;
        RECT 80.610 66.260 80.940 66.275 ;
        RECT 85.945 66.260 86.275 66.275 ;
        RECT 91.270 66.260 91.600 66.275 ;
        RECT 101.930 66.260 102.260 66.275 ;
        RECT 107.265 66.260 107.595 66.275 ;
        RECT 112.590 66.260 112.920 66.275 ;
        RECT 117.925 66.260 118.255 66.275 ;
        RECT 80.610 65.960 92.040 66.260 ;
        RECT 101.930 65.960 113.360 66.260 ;
        RECT 117.485 65.960 118.255 66.260 ;
        RECT 80.610 65.945 80.940 65.960 ;
        RECT 85.945 65.945 86.275 65.960 ;
        RECT 91.270 65.945 91.600 65.960 ;
        RECT 101.930 65.945 102.260 65.960 ;
        RECT 107.265 65.945 107.595 65.960 ;
        RECT 112.590 65.945 112.920 65.960 ;
        RECT 117.925 65.945 118.255 65.960 ;
        RECT 29.735 65.555 30.935 65.570 ;
        RECT 31.480 65.555 31.810 65.570 ;
        RECT 36.805 65.555 37.135 65.570 ;
        RECT 42.140 65.555 42.470 65.570 ;
        RECT 47.465 65.555 47.795 65.570 ;
        RECT 52.800 65.555 53.130 65.570 ;
        RECT 58.125 65.555 58.455 65.570 ;
        RECT 63.460 65.555 63.790 65.570 ;
        RECT 68.785 65.555 69.115 65.570 ;
        RECT 74.120 65.555 74.450 65.570 ;
        RECT 79.445 65.555 79.775 65.570 ;
        RECT 84.780 65.555 85.110 65.570 ;
        RECT 90.105 65.555 90.435 65.570 ;
        RECT 95.440 65.555 95.770 65.570 ;
        RECT 100.765 65.555 101.095 65.570 ;
        RECT 106.100 65.555 106.430 65.570 ;
        RECT 111.425 65.555 111.755 65.570 ;
        RECT 116.760 65.555 117.090 65.570 ;
        RECT 122.085 65.555 122.415 65.570 ;
        RECT 29.705 65.255 127.180 65.555 ;
        RECT 29.735 65.240 30.935 65.255 ;
        RECT 31.480 65.240 31.810 65.255 ;
        RECT 36.805 65.240 37.135 65.255 ;
        RECT 42.140 65.240 42.470 65.255 ;
        RECT 47.465 65.240 47.795 65.255 ;
        RECT 52.800 65.240 53.130 65.255 ;
        RECT 58.125 65.240 58.455 65.255 ;
        RECT 63.460 65.240 63.790 65.255 ;
        RECT 68.785 65.240 69.115 65.255 ;
        RECT 74.120 65.240 74.450 65.255 ;
        RECT 79.445 65.240 79.775 65.255 ;
        RECT 84.780 65.240 85.110 65.255 ;
        RECT 90.105 65.240 90.435 65.255 ;
        RECT 95.440 65.240 95.770 65.255 ;
        RECT 100.765 65.240 101.095 65.255 ;
        RECT 106.100 65.240 106.430 65.255 ;
        RECT 111.425 65.240 111.755 65.255 ;
        RECT 116.760 65.240 117.090 65.255 ;
        RECT 122.085 65.240 122.415 65.255 ;
        RECT 29.735 64.910 30.935 64.925 ;
        RECT 35.980 64.910 36.310 64.925 ;
        RECT 41.305 64.910 41.635 64.925 ;
        RECT 46.640 64.910 46.970 64.925 ;
        RECT 51.965 64.910 52.295 64.925 ;
        RECT 57.300 64.910 57.630 64.925 ;
        RECT 62.625 64.910 62.955 64.925 ;
        RECT 67.960 64.910 68.290 64.925 ;
        RECT 73.285 64.910 73.615 64.925 ;
        RECT 78.620 64.910 78.950 64.925 ;
        RECT 83.945 64.910 84.275 64.925 ;
        RECT 89.280 64.910 89.610 64.925 ;
        RECT 94.605 64.910 94.935 64.925 ;
        RECT 99.940 64.910 100.270 64.925 ;
        RECT 105.265 64.910 105.595 64.925 ;
        RECT 110.600 64.910 110.930 64.925 ;
        RECT 115.925 64.910 116.255 64.925 ;
        RECT 121.260 64.910 121.590 64.925 ;
        RECT 126.585 64.910 126.915 64.925 ;
        RECT 29.705 64.610 127.180 64.910 ;
        RECT 29.735 64.595 30.935 64.610 ;
        RECT 35.980 64.595 36.310 64.610 ;
        RECT 41.305 64.595 41.635 64.610 ;
        RECT 46.640 64.595 46.970 64.610 ;
        RECT 51.965 64.595 52.295 64.610 ;
        RECT 57.300 64.595 57.630 64.610 ;
        RECT 62.625 64.595 62.955 64.610 ;
        RECT 67.960 64.595 68.290 64.610 ;
        RECT 73.285 64.595 73.615 64.610 ;
        RECT 78.620 64.595 78.950 64.610 ;
        RECT 83.945 64.595 84.275 64.610 ;
        RECT 89.280 64.595 89.610 64.610 ;
        RECT 94.605 64.595 94.935 64.610 ;
        RECT 99.940 64.595 100.270 64.610 ;
        RECT 105.265 64.595 105.595 64.610 ;
        RECT 110.600 64.595 110.930 64.610 ;
        RECT 115.925 64.595 116.255 64.610 ;
        RECT 121.260 64.595 121.590 64.610 ;
        RECT 126.585 64.595 126.915 64.610 ;
        RECT 29.735 64.265 30.935 64.280 ;
        RECT 31.480 64.265 31.810 64.275 ;
        RECT 36.805 64.265 37.135 64.275 ;
        RECT 42.140 64.265 42.470 64.275 ;
        RECT 47.465 64.265 47.795 64.275 ;
        RECT 52.800 64.265 53.130 64.275 ;
        RECT 58.125 64.265 58.455 64.275 ;
        RECT 63.460 64.265 63.790 64.275 ;
        RECT 68.785 64.265 69.115 64.275 ;
        RECT 74.120 64.265 74.450 64.275 ;
        RECT 79.445 64.265 79.775 64.275 ;
        RECT 84.780 64.265 85.110 64.275 ;
        RECT 90.105 64.265 90.435 64.275 ;
        RECT 95.440 64.265 95.770 64.275 ;
        RECT 100.765 64.265 101.095 64.275 ;
        RECT 106.100 64.265 106.430 64.275 ;
        RECT 111.425 64.265 111.755 64.275 ;
        RECT 116.760 64.265 117.090 64.275 ;
        RECT 122.085 64.265 122.415 64.275 ;
        RECT 29.705 63.965 127.180 64.265 ;
        RECT 29.735 63.950 30.935 63.965 ;
        RECT 31.480 63.945 31.810 63.965 ;
        RECT 36.805 63.945 37.135 63.965 ;
        RECT 42.140 63.945 42.470 63.965 ;
        RECT 47.465 63.945 47.795 63.965 ;
        RECT 52.800 63.945 53.130 63.965 ;
        RECT 58.125 63.945 58.455 63.965 ;
        RECT 63.460 63.945 63.790 63.965 ;
        RECT 68.785 63.945 69.115 63.965 ;
        RECT 74.120 63.945 74.450 63.965 ;
        RECT 79.445 63.945 79.775 63.965 ;
        RECT 84.780 63.945 85.110 63.965 ;
        RECT 90.105 63.945 90.435 63.965 ;
        RECT 95.440 63.945 95.770 63.965 ;
        RECT 100.765 63.945 101.095 63.965 ;
        RECT 106.100 63.945 106.430 63.965 ;
        RECT 111.425 63.945 111.755 63.965 ;
        RECT 116.760 63.945 117.090 63.965 ;
        RECT 122.085 63.945 122.415 63.965 ;
        RECT 29.735 63.620 30.935 63.635 ;
        RECT 35.985 63.620 36.315 63.645 ;
        RECT 41.310 63.620 41.640 63.645 ;
        RECT 46.645 63.620 46.975 63.645 ;
        RECT 51.970 63.620 52.300 63.645 ;
        RECT 57.305 63.620 57.635 63.645 ;
        RECT 62.630 63.620 62.960 63.645 ;
        RECT 67.965 63.620 68.295 63.645 ;
        RECT 73.290 63.620 73.620 63.645 ;
        RECT 78.625 63.620 78.955 63.645 ;
        RECT 83.950 63.620 84.280 63.645 ;
        RECT 89.285 63.620 89.615 63.645 ;
        RECT 94.610 63.620 94.940 63.645 ;
        RECT 99.945 63.620 100.275 63.645 ;
        RECT 105.270 63.620 105.600 63.645 ;
        RECT 110.605 63.620 110.935 63.645 ;
        RECT 115.930 63.620 116.260 63.645 ;
        RECT 121.265 63.620 121.595 63.645 ;
        RECT 126.590 63.620 126.920 63.645 ;
        RECT 29.705 63.320 127.180 63.620 ;
        RECT 29.735 63.305 30.935 63.320 ;
        RECT 35.985 63.315 36.315 63.320 ;
        RECT 41.310 63.315 41.640 63.320 ;
        RECT 46.645 63.315 46.975 63.320 ;
        RECT 51.970 63.315 52.300 63.320 ;
        RECT 57.305 63.315 57.635 63.320 ;
        RECT 62.630 63.315 62.960 63.320 ;
        RECT 67.965 63.315 68.295 63.320 ;
        RECT 73.290 63.315 73.620 63.320 ;
        RECT 78.625 63.315 78.955 63.320 ;
        RECT 83.950 63.315 84.280 63.320 ;
        RECT 89.285 63.315 89.615 63.320 ;
        RECT 94.610 63.315 94.940 63.320 ;
        RECT 99.945 63.315 100.275 63.320 ;
        RECT 105.270 63.315 105.600 63.320 ;
        RECT 110.605 63.315 110.935 63.320 ;
        RECT 115.930 63.315 116.260 63.320 ;
        RECT 121.265 63.315 121.595 63.320 ;
        RECT 126.590 63.315 126.920 63.320 ;
        RECT 29.735 61.290 30.935 61.305 ;
        RECT 31.485 61.290 31.815 61.305 ;
        RECT 36.810 61.290 37.140 61.305 ;
        RECT 42.145 61.290 42.475 61.305 ;
        RECT 47.470 61.290 47.800 61.305 ;
        RECT 52.805 61.290 53.135 61.305 ;
        RECT 58.130 61.290 58.460 61.305 ;
        RECT 63.465 61.290 63.795 61.305 ;
        RECT 68.790 61.290 69.120 61.305 ;
        RECT 74.125 61.290 74.455 61.305 ;
        RECT 79.450 61.290 79.780 61.305 ;
        RECT 84.785 61.290 85.115 61.305 ;
        RECT 90.110 61.290 90.440 61.305 ;
        RECT 95.445 61.290 95.775 61.305 ;
        RECT 100.770 61.290 101.100 61.305 ;
        RECT 106.105 61.290 106.435 61.305 ;
        RECT 111.430 61.290 111.760 61.305 ;
        RECT 116.765 61.290 117.095 61.305 ;
        RECT 122.090 61.290 122.420 61.305 ;
        RECT 29.705 60.990 127.180 61.290 ;
        RECT 29.735 60.975 30.935 60.990 ;
        RECT 31.485 60.975 31.815 60.990 ;
        RECT 36.810 60.975 37.140 60.990 ;
        RECT 42.145 60.975 42.475 60.990 ;
        RECT 47.470 60.975 47.800 60.990 ;
        RECT 52.805 60.975 53.135 60.990 ;
        RECT 58.130 60.975 58.460 60.990 ;
        RECT 63.465 60.975 63.795 60.990 ;
        RECT 68.790 60.975 69.120 60.990 ;
        RECT 74.125 60.975 74.455 60.990 ;
        RECT 79.450 60.975 79.780 60.990 ;
        RECT 84.785 60.975 85.115 60.990 ;
        RECT 90.110 60.975 90.440 60.990 ;
        RECT 95.445 60.975 95.775 60.990 ;
        RECT 100.770 60.975 101.100 60.990 ;
        RECT 106.105 60.975 106.435 60.990 ;
        RECT 111.430 60.975 111.760 60.990 ;
        RECT 116.765 60.975 117.095 60.990 ;
        RECT 122.090 60.975 122.420 60.990 ;
        RECT 29.735 60.645 30.935 60.660 ;
        RECT 35.980 60.645 36.310 60.660 ;
        RECT 41.305 60.645 41.635 60.660 ;
        RECT 46.640 60.645 46.970 60.660 ;
        RECT 51.965 60.645 52.295 60.660 ;
        RECT 57.300 60.645 57.630 60.660 ;
        RECT 62.625 60.645 62.955 60.660 ;
        RECT 67.960 60.645 68.290 60.660 ;
        RECT 73.285 60.645 73.615 60.660 ;
        RECT 78.620 60.645 78.950 60.660 ;
        RECT 83.945 60.645 84.275 60.660 ;
        RECT 89.280 60.645 89.610 60.660 ;
        RECT 94.605 60.645 94.935 60.660 ;
        RECT 99.940 60.645 100.270 60.660 ;
        RECT 105.265 60.645 105.595 60.660 ;
        RECT 110.600 60.645 110.930 60.660 ;
        RECT 115.925 60.645 116.255 60.660 ;
        RECT 121.260 60.645 121.590 60.660 ;
        RECT 126.585 60.645 126.915 60.660 ;
        RECT 29.705 60.345 127.180 60.645 ;
        RECT 29.735 60.330 30.935 60.345 ;
        RECT 35.980 60.330 36.310 60.345 ;
        RECT 41.305 60.330 41.635 60.345 ;
        RECT 46.640 60.330 46.970 60.345 ;
        RECT 51.965 60.330 52.295 60.345 ;
        RECT 57.300 60.330 57.630 60.345 ;
        RECT 62.625 60.330 62.955 60.345 ;
        RECT 67.960 60.330 68.290 60.345 ;
        RECT 73.285 60.330 73.615 60.345 ;
        RECT 78.620 60.330 78.950 60.345 ;
        RECT 83.945 60.330 84.275 60.345 ;
        RECT 89.280 60.330 89.610 60.345 ;
        RECT 94.605 60.330 94.935 60.345 ;
        RECT 99.940 60.330 100.270 60.345 ;
        RECT 105.265 60.330 105.595 60.345 ;
        RECT 110.600 60.330 110.930 60.345 ;
        RECT 115.925 60.330 116.255 60.345 ;
        RECT 121.260 60.330 121.590 60.345 ;
        RECT 126.585 60.330 126.915 60.345 ;
        RECT 29.735 60.000 30.935 60.015 ;
        RECT 31.480 60.000 31.810 60.015 ;
        RECT 36.805 60.000 37.135 60.015 ;
        RECT 42.140 60.000 42.470 60.015 ;
        RECT 47.465 60.000 47.795 60.015 ;
        RECT 52.800 60.000 53.130 60.015 ;
        RECT 58.125 60.000 58.455 60.015 ;
        RECT 63.460 60.000 63.790 60.015 ;
        RECT 68.785 60.000 69.115 60.015 ;
        RECT 74.120 60.000 74.450 60.015 ;
        RECT 79.445 60.000 79.775 60.015 ;
        RECT 84.780 60.000 85.110 60.015 ;
        RECT 90.105 60.000 90.435 60.015 ;
        RECT 95.440 60.000 95.770 60.015 ;
        RECT 100.765 60.000 101.095 60.015 ;
        RECT 106.100 60.000 106.430 60.015 ;
        RECT 111.425 60.000 111.755 60.015 ;
        RECT 116.760 60.000 117.090 60.015 ;
        RECT 122.085 60.000 122.415 60.015 ;
        RECT 29.705 59.700 127.180 60.000 ;
        RECT 29.735 59.685 30.935 59.700 ;
        RECT 31.480 59.685 31.810 59.700 ;
        RECT 36.805 59.685 37.135 59.700 ;
        RECT 42.140 59.685 42.470 59.700 ;
        RECT 47.465 59.685 47.795 59.700 ;
        RECT 52.800 59.685 53.130 59.700 ;
        RECT 58.125 59.685 58.455 59.700 ;
        RECT 63.460 59.685 63.790 59.700 ;
        RECT 68.785 59.685 69.115 59.700 ;
        RECT 74.120 59.685 74.450 59.700 ;
        RECT 79.445 59.685 79.775 59.700 ;
        RECT 84.780 59.685 85.110 59.700 ;
        RECT 90.105 59.685 90.435 59.700 ;
        RECT 95.440 59.685 95.770 59.700 ;
        RECT 100.765 59.685 101.095 59.700 ;
        RECT 106.100 59.685 106.430 59.700 ;
        RECT 111.425 59.685 111.755 59.700 ;
        RECT 116.760 59.685 117.090 59.700 ;
        RECT 122.085 59.685 122.415 59.700 ;
        RECT 29.735 59.355 30.935 59.370 ;
        RECT 35.980 59.355 36.310 59.370 ;
        RECT 41.305 59.355 41.635 59.370 ;
        RECT 46.640 59.355 46.970 59.370 ;
        RECT 51.965 59.355 52.295 59.370 ;
        RECT 57.300 59.355 57.630 59.370 ;
        RECT 62.625 59.355 62.955 59.370 ;
        RECT 67.960 59.355 68.290 59.370 ;
        RECT 73.285 59.355 73.615 59.370 ;
        RECT 78.620 59.355 78.950 59.370 ;
        RECT 83.945 59.355 84.275 59.370 ;
        RECT 89.280 59.355 89.610 59.370 ;
        RECT 94.605 59.355 94.935 59.370 ;
        RECT 99.940 59.355 100.270 59.370 ;
        RECT 105.265 59.355 105.595 59.370 ;
        RECT 110.600 59.355 110.930 59.370 ;
        RECT 115.925 59.355 116.255 59.370 ;
        RECT 121.260 59.355 121.590 59.370 ;
        RECT 126.585 59.355 126.915 59.370 ;
        RECT 29.705 59.055 127.180 59.355 ;
        RECT 29.735 59.040 30.935 59.055 ;
        RECT 35.980 59.040 36.310 59.055 ;
        RECT 41.305 59.040 41.635 59.055 ;
        RECT 46.640 59.040 46.970 59.055 ;
        RECT 51.965 59.040 52.295 59.055 ;
        RECT 57.300 59.040 57.630 59.055 ;
        RECT 62.625 59.040 62.955 59.055 ;
        RECT 67.960 59.040 68.290 59.055 ;
        RECT 73.285 59.040 73.615 59.055 ;
        RECT 78.620 59.040 78.950 59.055 ;
        RECT 83.945 59.040 84.275 59.055 ;
        RECT 89.280 59.040 89.610 59.055 ;
        RECT 94.605 59.040 94.935 59.055 ;
        RECT 99.940 59.040 100.270 59.055 ;
        RECT 105.265 59.040 105.595 59.055 ;
        RECT 110.600 59.040 110.930 59.055 ;
        RECT 115.925 59.040 116.255 59.055 ;
        RECT 121.260 59.040 121.590 59.055 ;
        RECT 126.585 59.040 126.915 59.055 ;
        RECT 29.735 58.020 30.935 58.035 ;
        RECT 31.480 58.020 31.810 58.035 ;
        RECT 36.805 58.020 37.135 58.035 ;
        RECT 42.140 58.020 42.470 58.035 ;
        RECT 47.465 58.020 47.795 58.035 ;
        RECT 52.800 58.020 53.130 58.035 ;
        RECT 58.125 58.020 58.455 58.035 ;
        RECT 63.460 58.020 63.790 58.035 ;
        RECT 68.785 58.020 69.115 58.035 ;
        RECT 74.120 58.020 74.450 58.035 ;
        RECT 79.445 58.020 79.775 58.035 ;
        RECT 84.780 58.020 85.110 58.035 ;
        RECT 90.105 58.020 90.435 58.035 ;
        RECT 95.440 58.020 95.770 58.035 ;
        RECT 100.765 58.020 101.095 58.035 ;
        RECT 106.100 58.020 106.430 58.035 ;
        RECT 111.425 58.020 111.755 58.035 ;
        RECT 116.760 58.020 117.090 58.035 ;
        RECT 122.085 58.020 122.415 58.035 ;
        RECT 29.705 57.720 127.180 58.020 ;
        RECT 29.735 57.705 30.935 57.720 ;
        RECT 31.480 57.705 31.810 57.720 ;
        RECT 36.805 57.705 37.135 57.720 ;
        RECT 42.140 57.705 42.470 57.720 ;
        RECT 47.465 57.705 47.795 57.720 ;
        RECT 52.800 57.705 53.130 57.720 ;
        RECT 58.125 57.705 58.455 57.720 ;
        RECT 63.460 57.705 63.790 57.720 ;
        RECT 68.785 57.705 69.115 57.720 ;
        RECT 74.120 57.705 74.450 57.720 ;
        RECT 79.445 57.705 79.775 57.720 ;
        RECT 84.780 57.705 85.110 57.720 ;
        RECT 90.105 57.705 90.435 57.720 ;
        RECT 95.440 57.705 95.770 57.720 ;
        RECT 100.765 57.705 101.095 57.720 ;
        RECT 106.100 57.705 106.430 57.720 ;
        RECT 111.425 57.705 111.755 57.720 ;
        RECT 116.760 57.705 117.090 57.720 ;
        RECT 122.085 57.705 122.415 57.720 ;
        RECT 29.735 57.375 30.935 57.390 ;
        RECT 35.980 57.375 36.310 57.390 ;
        RECT 41.305 57.375 41.635 57.390 ;
        RECT 46.640 57.375 46.970 57.390 ;
        RECT 51.965 57.375 52.295 57.390 ;
        RECT 57.300 57.375 57.630 57.390 ;
        RECT 62.625 57.375 62.955 57.390 ;
        RECT 67.960 57.375 68.290 57.390 ;
        RECT 73.285 57.375 73.615 57.390 ;
        RECT 78.620 57.375 78.950 57.390 ;
        RECT 83.945 57.375 84.275 57.390 ;
        RECT 89.280 57.375 89.610 57.390 ;
        RECT 94.605 57.375 94.935 57.390 ;
        RECT 99.940 57.375 100.270 57.390 ;
        RECT 105.265 57.375 105.595 57.390 ;
        RECT 110.600 57.375 110.930 57.390 ;
        RECT 115.925 57.375 116.255 57.390 ;
        RECT 121.260 57.375 121.590 57.390 ;
        RECT 126.585 57.375 126.915 57.390 ;
        RECT 29.705 57.075 127.180 57.375 ;
        RECT 29.735 57.060 30.935 57.075 ;
        RECT 35.980 57.060 36.310 57.075 ;
        RECT 41.305 57.060 41.635 57.075 ;
        RECT 46.640 57.060 46.970 57.075 ;
        RECT 51.965 57.060 52.295 57.075 ;
        RECT 57.300 57.060 57.630 57.075 ;
        RECT 62.625 57.060 62.955 57.075 ;
        RECT 67.960 57.060 68.290 57.075 ;
        RECT 73.285 57.060 73.615 57.075 ;
        RECT 78.620 57.060 78.950 57.075 ;
        RECT 83.945 57.060 84.275 57.075 ;
        RECT 89.280 57.060 89.610 57.075 ;
        RECT 94.605 57.060 94.935 57.075 ;
        RECT 99.940 57.060 100.270 57.075 ;
        RECT 105.265 57.060 105.595 57.075 ;
        RECT 110.600 57.060 110.930 57.075 ;
        RECT 115.925 57.060 116.255 57.075 ;
        RECT 121.260 57.060 121.590 57.075 ;
        RECT 126.585 57.060 126.915 57.075 ;
        RECT 29.735 56.730 30.935 56.745 ;
        RECT 31.480 56.730 31.810 56.740 ;
        RECT 36.805 56.730 37.135 56.740 ;
        RECT 42.140 56.730 42.470 56.740 ;
        RECT 47.465 56.730 47.795 56.740 ;
        RECT 52.800 56.730 53.130 56.740 ;
        RECT 58.125 56.730 58.455 56.740 ;
        RECT 63.460 56.730 63.790 56.740 ;
        RECT 68.785 56.730 69.115 56.740 ;
        RECT 74.120 56.730 74.450 56.740 ;
        RECT 79.445 56.730 79.775 56.740 ;
        RECT 84.780 56.730 85.110 56.740 ;
        RECT 90.105 56.730 90.435 56.740 ;
        RECT 95.440 56.730 95.770 56.740 ;
        RECT 100.765 56.730 101.095 56.740 ;
        RECT 106.100 56.730 106.430 56.740 ;
        RECT 111.425 56.730 111.755 56.740 ;
        RECT 116.760 56.730 117.090 56.740 ;
        RECT 122.085 56.730 122.415 56.740 ;
        RECT 29.705 56.430 127.180 56.730 ;
        RECT 29.735 56.415 30.935 56.430 ;
        RECT 31.480 56.410 31.810 56.430 ;
        RECT 36.805 56.410 37.135 56.430 ;
        RECT 42.140 56.410 42.470 56.430 ;
        RECT 47.465 56.410 47.795 56.430 ;
        RECT 52.800 56.410 53.130 56.430 ;
        RECT 58.125 56.410 58.455 56.430 ;
        RECT 63.460 56.410 63.790 56.430 ;
        RECT 68.785 56.410 69.115 56.430 ;
        RECT 74.120 56.410 74.450 56.430 ;
        RECT 79.445 56.410 79.775 56.430 ;
        RECT 84.780 56.410 85.110 56.430 ;
        RECT 90.105 56.410 90.435 56.430 ;
        RECT 95.440 56.410 95.770 56.430 ;
        RECT 100.765 56.410 101.095 56.430 ;
        RECT 106.100 56.410 106.430 56.430 ;
        RECT 111.425 56.410 111.755 56.430 ;
        RECT 116.760 56.410 117.090 56.430 ;
        RECT 122.085 56.410 122.415 56.430 ;
        RECT 29.735 56.085 30.935 56.100 ;
        RECT 35.985 56.085 36.315 56.110 ;
        RECT 41.310 56.085 41.640 56.110 ;
        RECT 46.645 56.085 46.975 56.110 ;
        RECT 51.970 56.085 52.300 56.110 ;
        RECT 57.305 56.085 57.635 56.110 ;
        RECT 62.630 56.085 62.960 56.110 ;
        RECT 67.965 56.085 68.295 56.110 ;
        RECT 73.290 56.085 73.620 56.110 ;
        RECT 78.625 56.085 78.955 56.110 ;
        RECT 83.950 56.085 84.280 56.110 ;
        RECT 89.285 56.085 89.615 56.110 ;
        RECT 94.610 56.085 94.940 56.110 ;
        RECT 99.945 56.085 100.275 56.110 ;
        RECT 105.270 56.085 105.600 56.110 ;
        RECT 110.605 56.085 110.935 56.110 ;
        RECT 115.930 56.085 116.260 56.110 ;
        RECT 121.265 56.085 121.595 56.110 ;
        RECT 126.590 56.085 126.920 56.110 ;
        RECT 29.705 55.785 127.180 56.085 ;
        RECT 29.735 55.770 30.935 55.785 ;
        RECT 35.985 55.780 36.315 55.785 ;
        RECT 41.310 55.780 41.640 55.785 ;
        RECT 46.645 55.780 46.975 55.785 ;
        RECT 51.970 55.780 52.300 55.785 ;
        RECT 57.305 55.780 57.635 55.785 ;
        RECT 62.630 55.780 62.960 55.785 ;
        RECT 67.965 55.780 68.295 55.785 ;
        RECT 73.290 55.780 73.620 55.785 ;
        RECT 78.625 55.780 78.955 55.785 ;
        RECT 83.950 55.780 84.280 55.785 ;
        RECT 89.285 55.780 89.615 55.785 ;
        RECT 94.610 55.780 94.940 55.785 ;
        RECT 99.945 55.780 100.275 55.785 ;
        RECT 105.270 55.780 105.600 55.785 ;
        RECT 110.605 55.780 110.935 55.785 ;
        RECT 115.930 55.780 116.260 55.785 ;
        RECT 121.265 55.780 121.595 55.785 ;
        RECT 126.590 55.780 126.920 55.785 ;
        RECT 29.735 53.755 30.935 53.770 ;
        RECT 31.485 53.755 31.815 53.770 ;
        RECT 36.810 53.755 37.140 53.770 ;
        RECT 42.145 53.755 42.475 53.770 ;
        RECT 47.470 53.755 47.800 53.770 ;
        RECT 52.805 53.755 53.135 53.770 ;
        RECT 58.130 53.755 58.460 53.770 ;
        RECT 63.465 53.755 63.795 53.770 ;
        RECT 68.790 53.755 69.120 53.770 ;
        RECT 74.125 53.755 74.455 53.770 ;
        RECT 79.450 53.755 79.780 53.770 ;
        RECT 84.785 53.755 85.115 53.770 ;
        RECT 90.110 53.755 90.440 53.770 ;
        RECT 95.445 53.755 95.775 53.770 ;
        RECT 100.770 53.755 101.100 53.770 ;
        RECT 106.105 53.755 106.435 53.770 ;
        RECT 111.430 53.755 111.760 53.770 ;
        RECT 116.765 53.755 117.095 53.770 ;
        RECT 122.090 53.755 122.420 53.770 ;
        RECT 29.705 53.455 127.180 53.755 ;
        RECT 29.735 53.440 30.935 53.455 ;
        RECT 31.485 53.440 31.815 53.455 ;
        RECT 36.810 53.440 37.140 53.455 ;
        RECT 42.145 53.440 42.475 53.455 ;
        RECT 47.470 53.440 47.800 53.455 ;
        RECT 52.805 53.440 53.135 53.455 ;
        RECT 58.130 53.440 58.460 53.455 ;
        RECT 63.465 53.440 63.795 53.455 ;
        RECT 68.790 53.440 69.120 53.455 ;
        RECT 74.125 53.440 74.455 53.455 ;
        RECT 79.450 53.440 79.780 53.455 ;
        RECT 84.785 53.440 85.115 53.455 ;
        RECT 90.110 53.440 90.440 53.455 ;
        RECT 95.445 53.440 95.775 53.455 ;
        RECT 100.770 53.440 101.100 53.455 ;
        RECT 106.105 53.440 106.435 53.455 ;
        RECT 111.430 53.440 111.760 53.455 ;
        RECT 116.765 53.440 117.095 53.455 ;
        RECT 122.090 53.440 122.420 53.455 ;
        RECT 29.735 53.110 30.935 53.125 ;
        RECT 35.980 53.110 36.310 53.125 ;
        RECT 41.305 53.110 41.635 53.125 ;
        RECT 46.640 53.110 46.970 53.125 ;
        RECT 51.965 53.110 52.295 53.125 ;
        RECT 57.300 53.110 57.630 53.125 ;
        RECT 62.625 53.110 62.955 53.125 ;
        RECT 67.960 53.110 68.290 53.125 ;
        RECT 73.285 53.110 73.615 53.125 ;
        RECT 78.620 53.110 78.950 53.125 ;
        RECT 83.945 53.110 84.275 53.125 ;
        RECT 89.280 53.110 89.610 53.125 ;
        RECT 94.605 53.110 94.935 53.125 ;
        RECT 99.940 53.110 100.270 53.125 ;
        RECT 105.265 53.110 105.595 53.125 ;
        RECT 110.600 53.110 110.930 53.125 ;
        RECT 115.925 53.110 116.255 53.125 ;
        RECT 121.260 53.110 121.590 53.125 ;
        RECT 126.585 53.110 126.915 53.125 ;
        RECT 29.705 52.810 127.180 53.110 ;
        RECT 29.735 52.795 30.935 52.810 ;
        RECT 35.980 52.795 36.310 52.810 ;
        RECT 41.305 52.795 41.635 52.810 ;
        RECT 46.640 52.795 46.970 52.810 ;
        RECT 51.965 52.795 52.295 52.810 ;
        RECT 57.300 52.795 57.630 52.810 ;
        RECT 62.625 52.795 62.955 52.810 ;
        RECT 67.960 52.795 68.290 52.810 ;
        RECT 73.285 52.795 73.615 52.810 ;
        RECT 78.620 52.795 78.950 52.810 ;
        RECT 83.945 52.795 84.275 52.810 ;
        RECT 89.280 52.795 89.610 52.810 ;
        RECT 94.605 52.795 94.935 52.810 ;
        RECT 99.940 52.795 100.270 52.810 ;
        RECT 105.265 52.795 105.595 52.810 ;
        RECT 110.600 52.795 110.930 52.810 ;
        RECT 115.925 52.795 116.255 52.810 ;
        RECT 121.260 52.795 121.590 52.810 ;
        RECT 126.585 52.795 126.915 52.810 ;
        RECT 29.735 52.465 30.935 52.480 ;
        RECT 31.480 52.465 31.810 52.480 ;
        RECT 36.805 52.465 37.135 52.480 ;
        RECT 42.140 52.465 42.470 52.480 ;
        RECT 47.465 52.465 47.795 52.480 ;
        RECT 52.800 52.465 53.130 52.480 ;
        RECT 58.125 52.465 58.455 52.480 ;
        RECT 63.460 52.465 63.790 52.480 ;
        RECT 68.785 52.465 69.115 52.480 ;
        RECT 74.120 52.465 74.450 52.480 ;
        RECT 79.445 52.465 79.775 52.480 ;
        RECT 84.780 52.465 85.110 52.480 ;
        RECT 90.105 52.465 90.435 52.480 ;
        RECT 95.440 52.465 95.770 52.480 ;
        RECT 100.765 52.465 101.095 52.480 ;
        RECT 106.100 52.465 106.430 52.480 ;
        RECT 111.425 52.465 111.755 52.480 ;
        RECT 116.760 52.465 117.090 52.480 ;
        RECT 122.085 52.465 122.415 52.480 ;
        RECT 29.705 52.165 127.180 52.465 ;
        RECT 29.735 52.150 30.935 52.165 ;
        RECT 31.480 52.150 31.810 52.165 ;
        RECT 36.805 52.150 37.135 52.165 ;
        RECT 42.140 52.150 42.470 52.165 ;
        RECT 47.465 52.150 47.795 52.165 ;
        RECT 52.800 52.150 53.130 52.165 ;
        RECT 58.125 52.150 58.455 52.165 ;
        RECT 63.460 52.150 63.790 52.165 ;
        RECT 68.785 52.150 69.115 52.165 ;
        RECT 74.120 52.150 74.450 52.165 ;
        RECT 79.445 52.150 79.775 52.165 ;
        RECT 84.780 52.150 85.110 52.165 ;
        RECT 90.105 52.150 90.435 52.165 ;
        RECT 95.440 52.150 95.770 52.165 ;
        RECT 100.765 52.150 101.095 52.165 ;
        RECT 106.100 52.150 106.430 52.165 ;
        RECT 111.425 52.150 111.755 52.165 ;
        RECT 116.760 52.150 117.090 52.165 ;
        RECT 122.085 52.150 122.415 52.165 ;
        RECT 29.735 51.820 30.935 51.835 ;
        RECT 35.980 51.820 36.310 51.835 ;
        RECT 41.305 51.820 41.635 51.835 ;
        RECT 46.640 51.820 46.970 51.835 ;
        RECT 51.965 51.820 52.295 51.835 ;
        RECT 57.300 51.820 57.630 51.835 ;
        RECT 62.625 51.820 62.955 51.835 ;
        RECT 67.960 51.820 68.290 51.835 ;
        RECT 73.285 51.820 73.615 51.835 ;
        RECT 78.620 51.820 78.950 51.835 ;
        RECT 83.945 51.820 84.275 51.835 ;
        RECT 89.280 51.820 89.610 51.835 ;
        RECT 94.605 51.820 94.935 51.835 ;
        RECT 99.940 51.820 100.270 51.835 ;
        RECT 105.265 51.820 105.595 51.835 ;
        RECT 110.600 51.820 110.930 51.835 ;
        RECT 115.925 51.820 116.255 51.835 ;
        RECT 121.260 51.820 121.590 51.835 ;
        RECT 126.585 51.820 126.915 51.835 ;
        RECT 29.705 51.520 127.180 51.820 ;
        RECT 29.735 51.505 30.935 51.520 ;
        RECT 35.980 51.505 36.310 51.520 ;
        RECT 41.305 51.505 41.635 51.520 ;
        RECT 46.640 51.505 46.970 51.520 ;
        RECT 51.965 51.505 52.295 51.520 ;
        RECT 57.300 51.505 57.630 51.520 ;
        RECT 62.625 51.505 62.955 51.520 ;
        RECT 67.960 51.505 68.290 51.520 ;
        RECT 73.285 51.505 73.615 51.520 ;
        RECT 78.620 51.505 78.950 51.520 ;
        RECT 83.945 51.505 84.275 51.520 ;
        RECT 89.280 51.505 89.610 51.520 ;
        RECT 94.605 51.505 94.935 51.520 ;
        RECT 99.940 51.505 100.270 51.520 ;
        RECT 105.265 51.505 105.595 51.520 ;
        RECT 110.600 51.505 110.930 51.520 ;
        RECT 115.925 51.505 116.255 51.520 ;
        RECT 121.260 51.505 121.590 51.520 ;
        RECT 126.585 51.505 126.915 51.520 ;
        RECT 29.735 50.485 30.935 50.500 ;
        RECT 31.480 50.485 31.810 50.500 ;
        RECT 36.805 50.485 37.135 50.500 ;
        RECT 42.140 50.485 42.470 50.500 ;
        RECT 47.465 50.485 47.795 50.500 ;
        RECT 52.800 50.485 53.130 50.500 ;
        RECT 58.125 50.485 58.455 50.500 ;
        RECT 63.460 50.485 63.790 50.500 ;
        RECT 68.785 50.485 69.115 50.500 ;
        RECT 74.120 50.485 74.450 50.500 ;
        RECT 79.445 50.485 79.775 50.500 ;
        RECT 84.780 50.485 85.110 50.500 ;
        RECT 90.105 50.485 90.435 50.500 ;
        RECT 95.440 50.485 95.770 50.500 ;
        RECT 100.765 50.485 101.095 50.500 ;
        RECT 106.100 50.485 106.430 50.500 ;
        RECT 111.425 50.485 111.755 50.500 ;
        RECT 116.760 50.485 117.090 50.500 ;
        RECT 122.085 50.485 122.415 50.500 ;
        RECT 29.705 50.185 127.180 50.485 ;
        RECT 29.735 50.170 30.935 50.185 ;
        RECT 31.480 50.170 31.810 50.185 ;
        RECT 36.805 50.170 37.135 50.185 ;
        RECT 42.140 50.170 42.470 50.185 ;
        RECT 47.465 50.170 47.795 50.185 ;
        RECT 52.800 50.170 53.130 50.185 ;
        RECT 58.125 50.170 58.455 50.185 ;
        RECT 63.460 50.170 63.790 50.185 ;
        RECT 68.785 50.170 69.115 50.185 ;
        RECT 74.120 50.170 74.450 50.185 ;
        RECT 79.445 50.170 79.775 50.185 ;
        RECT 84.780 50.170 85.110 50.185 ;
        RECT 90.105 50.170 90.435 50.185 ;
        RECT 95.440 50.170 95.770 50.185 ;
        RECT 100.765 50.170 101.095 50.185 ;
        RECT 106.100 50.170 106.430 50.185 ;
        RECT 111.425 50.170 111.755 50.185 ;
        RECT 116.760 50.170 117.090 50.185 ;
        RECT 122.085 50.170 122.415 50.185 ;
        RECT 29.735 49.840 30.935 49.855 ;
        RECT 35.980 49.840 36.310 49.855 ;
        RECT 41.305 49.840 41.635 49.855 ;
        RECT 46.640 49.840 46.970 49.855 ;
        RECT 51.965 49.840 52.295 49.855 ;
        RECT 57.300 49.840 57.630 49.855 ;
        RECT 62.625 49.840 62.955 49.855 ;
        RECT 67.960 49.840 68.290 49.855 ;
        RECT 73.285 49.840 73.615 49.855 ;
        RECT 78.620 49.840 78.950 49.855 ;
        RECT 83.945 49.840 84.275 49.855 ;
        RECT 89.280 49.840 89.610 49.855 ;
        RECT 94.605 49.840 94.935 49.855 ;
        RECT 99.940 49.840 100.270 49.855 ;
        RECT 105.265 49.840 105.595 49.855 ;
        RECT 110.600 49.840 110.930 49.855 ;
        RECT 115.925 49.840 116.255 49.855 ;
        RECT 121.260 49.840 121.590 49.855 ;
        RECT 126.585 49.840 126.915 49.855 ;
        RECT 29.705 49.540 127.180 49.840 ;
        RECT 29.735 49.525 30.935 49.540 ;
        RECT 35.980 49.525 36.310 49.540 ;
        RECT 41.305 49.525 41.635 49.540 ;
        RECT 46.640 49.525 46.970 49.540 ;
        RECT 51.965 49.525 52.295 49.540 ;
        RECT 57.300 49.525 57.630 49.540 ;
        RECT 62.625 49.525 62.955 49.540 ;
        RECT 67.960 49.525 68.290 49.540 ;
        RECT 73.285 49.525 73.615 49.540 ;
        RECT 78.620 49.525 78.950 49.540 ;
        RECT 83.945 49.525 84.275 49.540 ;
        RECT 89.280 49.525 89.610 49.540 ;
        RECT 94.605 49.525 94.935 49.540 ;
        RECT 99.940 49.525 100.270 49.540 ;
        RECT 105.265 49.525 105.595 49.540 ;
        RECT 110.600 49.525 110.930 49.540 ;
        RECT 115.925 49.525 116.255 49.540 ;
        RECT 121.260 49.525 121.590 49.540 ;
        RECT 126.585 49.525 126.915 49.540 ;
        RECT 29.735 49.195 30.935 49.210 ;
        RECT 31.480 49.195 31.810 49.205 ;
        RECT 36.805 49.195 37.135 49.205 ;
        RECT 42.140 49.195 42.470 49.205 ;
        RECT 47.465 49.195 47.795 49.205 ;
        RECT 52.800 49.195 53.130 49.205 ;
        RECT 58.125 49.195 58.455 49.205 ;
        RECT 63.460 49.195 63.790 49.205 ;
        RECT 68.785 49.195 69.115 49.205 ;
        RECT 74.120 49.195 74.450 49.205 ;
        RECT 79.445 49.195 79.775 49.205 ;
        RECT 84.780 49.195 85.110 49.205 ;
        RECT 90.105 49.195 90.435 49.205 ;
        RECT 95.440 49.195 95.770 49.205 ;
        RECT 100.765 49.195 101.095 49.205 ;
        RECT 106.100 49.195 106.430 49.205 ;
        RECT 111.425 49.195 111.755 49.205 ;
        RECT 116.760 49.195 117.090 49.205 ;
        RECT 122.085 49.195 122.415 49.205 ;
        RECT 29.705 48.895 127.180 49.195 ;
        RECT 29.735 48.880 30.935 48.895 ;
        RECT 31.480 48.875 31.810 48.895 ;
        RECT 36.805 48.875 37.135 48.895 ;
        RECT 42.140 48.875 42.470 48.895 ;
        RECT 47.465 48.875 47.795 48.895 ;
        RECT 52.800 48.875 53.130 48.895 ;
        RECT 58.125 48.875 58.455 48.895 ;
        RECT 63.460 48.875 63.790 48.895 ;
        RECT 68.785 48.875 69.115 48.895 ;
        RECT 74.120 48.875 74.450 48.895 ;
        RECT 79.445 48.875 79.775 48.895 ;
        RECT 84.780 48.875 85.110 48.895 ;
        RECT 90.105 48.875 90.435 48.895 ;
        RECT 95.440 48.875 95.770 48.895 ;
        RECT 100.765 48.875 101.095 48.895 ;
        RECT 106.100 48.875 106.430 48.895 ;
        RECT 111.425 48.875 111.755 48.895 ;
        RECT 116.760 48.875 117.090 48.895 ;
        RECT 122.085 48.875 122.415 48.895 ;
        RECT 29.735 48.550 30.935 48.565 ;
        RECT 35.985 48.550 36.315 48.575 ;
        RECT 41.310 48.550 41.640 48.575 ;
        RECT 46.645 48.550 46.975 48.575 ;
        RECT 51.970 48.550 52.300 48.575 ;
        RECT 57.305 48.550 57.635 48.575 ;
        RECT 62.630 48.550 62.960 48.575 ;
        RECT 67.965 48.550 68.295 48.575 ;
        RECT 73.290 48.550 73.620 48.575 ;
        RECT 78.625 48.550 78.955 48.575 ;
        RECT 83.950 48.550 84.280 48.575 ;
        RECT 89.285 48.550 89.615 48.575 ;
        RECT 94.610 48.550 94.940 48.575 ;
        RECT 99.945 48.550 100.275 48.575 ;
        RECT 105.270 48.550 105.600 48.575 ;
        RECT 110.605 48.550 110.935 48.575 ;
        RECT 115.930 48.550 116.260 48.575 ;
        RECT 121.265 48.550 121.595 48.575 ;
        RECT 126.590 48.550 126.920 48.575 ;
        RECT 29.705 48.250 127.180 48.550 ;
        RECT 29.735 48.235 30.935 48.250 ;
        RECT 35.985 48.245 36.315 48.250 ;
        RECT 41.310 48.245 41.640 48.250 ;
        RECT 46.645 48.245 46.975 48.250 ;
        RECT 51.970 48.245 52.300 48.250 ;
        RECT 57.305 48.245 57.635 48.250 ;
        RECT 62.630 48.245 62.960 48.250 ;
        RECT 67.965 48.245 68.295 48.250 ;
        RECT 73.290 48.245 73.620 48.250 ;
        RECT 78.625 48.245 78.955 48.250 ;
        RECT 83.950 48.245 84.280 48.250 ;
        RECT 89.285 48.245 89.615 48.250 ;
        RECT 94.610 48.245 94.940 48.250 ;
        RECT 99.945 48.245 100.275 48.250 ;
        RECT 105.270 48.245 105.600 48.250 ;
        RECT 110.605 48.245 110.935 48.250 ;
        RECT 115.930 48.245 116.260 48.250 ;
        RECT 121.265 48.245 121.595 48.250 ;
        RECT 126.590 48.245 126.920 48.250 ;
        RECT 29.735 46.220 30.935 46.235 ;
        RECT 31.485 46.220 31.815 46.235 ;
        RECT 36.810 46.220 37.140 46.235 ;
        RECT 42.145 46.220 42.475 46.235 ;
        RECT 47.470 46.220 47.800 46.235 ;
        RECT 52.805 46.220 53.135 46.235 ;
        RECT 58.130 46.220 58.460 46.235 ;
        RECT 63.465 46.220 63.795 46.235 ;
        RECT 68.790 46.220 69.120 46.235 ;
        RECT 74.125 46.220 74.455 46.235 ;
        RECT 79.450 46.220 79.780 46.235 ;
        RECT 84.785 46.220 85.115 46.235 ;
        RECT 90.110 46.220 90.440 46.235 ;
        RECT 95.445 46.220 95.775 46.235 ;
        RECT 100.770 46.220 101.100 46.235 ;
        RECT 106.105 46.220 106.435 46.235 ;
        RECT 111.430 46.220 111.760 46.235 ;
        RECT 116.765 46.220 117.095 46.235 ;
        RECT 122.090 46.220 122.420 46.235 ;
        RECT 29.705 45.920 127.180 46.220 ;
        RECT 29.735 45.905 30.935 45.920 ;
        RECT 31.485 45.905 31.815 45.920 ;
        RECT 36.810 45.905 37.140 45.920 ;
        RECT 42.145 45.905 42.475 45.920 ;
        RECT 47.470 45.905 47.800 45.920 ;
        RECT 52.805 45.905 53.135 45.920 ;
        RECT 58.130 45.905 58.460 45.920 ;
        RECT 63.465 45.905 63.795 45.920 ;
        RECT 68.790 45.905 69.120 45.920 ;
        RECT 74.125 45.905 74.455 45.920 ;
        RECT 79.450 45.905 79.780 45.920 ;
        RECT 84.785 45.905 85.115 45.920 ;
        RECT 90.110 45.905 90.440 45.920 ;
        RECT 95.445 45.905 95.775 45.920 ;
        RECT 100.770 45.905 101.100 45.920 ;
        RECT 106.105 45.905 106.435 45.920 ;
        RECT 111.430 45.905 111.760 45.920 ;
        RECT 116.765 45.905 117.095 45.920 ;
        RECT 122.090 45.905 122.420 45.920 ;
        RECT 29.735 45.575 30.935 45.590 ;
        RECT 35.980 45.575 36.310 45.590 ;
        RECT 41.305 45.575 41.635 45.590 ;
        RECT 46.640 45.575 46.970 45.590 ;
        RECT 51.965 45.575 52.295 45.590 ;
        RECT 57.300 45.575 57.630 45.590 ;
        RECT 62.625 45.575 62.955 45.590 ;
        RECT 67.960 45.575 68.290 45.590 ;
        RECT 73.285 45.575 73.615 45.590 ;
        RECT 78.620 45.575 78.950 45.590 ;
        RECT 83.945 45.575 84.275 45.590 ;
        RECT 89.280 45.575 89.610 45.590 ;
        RECT 94.605 45.575 94.935 45.590 ;
        RECT 99.940 45.575 100.270 45.590 ;
        RECT 105.265 45.575 105.595 45.590 ;
        RECT 110.600 45.575 110.930 45.590 ;
        RECT 115.925 45.575 116.255 45.590 ;
        RECT 121.260 45.575 121.590 45.590 ;
        RECT 126.585 45.575 126.915 45.590 ;
        RECT 29.705 45.275 127.180 45.575 ;
        RECT 29.735 45.260 30.935 45.275 ;
        RECT 35.980 45.260 36.310 45.275 ;
        RECT 41.305 45.260 41.635 45.275 ;
        RECT 46.640 45.260 46.970 45.275 ;
        RECT 51.965 45.260 52.295 45.275 ;
        RECT 57.300 45.260 57.630 45.275 ;
        RECT 62.625 45.260 62.955 45.275 ;
        RECT 67.960 45.260 68.290 45.275 ;
        RECT 73.285 45.260 73.615 45.275 ;
        RECT 78.620 45.260 78.950 45.275 ;
        RECT 83.945 45.260 84.275 45.275 ;
        RECT 89.280 45.260 89.610 45.275 ;
        RECT 94.605 45.260 94.935 45.275 ;
        RECT 99.940 45.260 100.270 45.275 ;
        RECT 105.265 45.260 105.595 45.275 ;
        RECT 110.600 45.260 110.930 45.275 ;
        RECT 115.925 45.260 116.255 45.275 ;
        RECT 121.260 45.260 121.590 45.275 ;
        RECT 126.585 45.260 126.915 45.275 ;
        RECT 29.735 44.930 30.935 44.945 ;
        RECT 31.480 44.930 31.810 44.945 ;
        RECT 36.805 44.930 37.135 44.945 ;
        RECT 42.140 44.930 42.470 44.945 ;
        RECT 47.465 44.930 47.795 44.945 ;
        RECT 52.800 44.930 53.130 44.945 ;
        RECT 58.125 44.930 58.455 44.945 ;
        RECT 63.460 44.930 63.790 44.945 ;
        RECT 68.785 44.930 69.115 44.945 ;
        RECT 74.120 44.930 74.450 44.945 ;
        RECT 79.445 44.930 79.775 44.945 ;
        RECT 84.780 44.930 85.110 44.945 ;
        RECT 90.105 44.930 90.435 44.945 ;
        RECT 95.440 44.930 95.770 44.945 ;
        RECT 100.765 44.930 101.095 44.945 ;
        RECT 106.100 44.930 106.430 44.945 ;
        RECT 111.425 44.930 111.755 44.945 ;
        RECT 116.760 44.930 117.090 44.945 ;
        RECT 122.085 44.930 122.415 44.945 ;
        RECT 29.705 44.630 127.180 44.930 ;
        RECT 29.735 44.615 30.935 44.630 ;
        RECT 31.480 44.615 31.810 44.630 ;
        RECT 36.805 44.615 37.135 44.630 ;
        RECT 42.140 44.615 42.470 44.630 ;
        RECT 47.465 44.615 47.795 44.630 ;
        RECT 52.800 44.615 53.130 44.630 ;
        RECT 58.125 44.615 58.455 44.630 ;
        RECT 63.460 44.615 63.790 44.630 ;
        RECT 68.785 44.615 69.115 44.630 ;
        RECT 74.120 44.615 74.450 44.630 ;
        RECT 79.445 44.615 79.775 44.630 ;
        RECT 84.780 44.615 85.110 44.630 ;
        RECT 90.105 44.615 90.435 44.630 ;
        RECT 95.440 44.615 95.770 44.630 ;
        RECT 100.765 44.615 101.095 44.630 ;
        RECT 106.100 44.615 106.430 44.630 ;
        RECT 111.425 44.615 111.755 44.630 ;
        RECT 116.760 44.615 117.090 44.630 ;
        RECT 122.085 44.615 122.415 44.630 ;
        RECT 29.735 44.285 30.935 44.300 ;
        RECT 35.980 44.285 36.310 44.300 ;
        RECT 41.305 44.285 41.635 44.300 ;
        RECT 46.640 44.285 46.970 44.300 ;
        RECT 51.965 44.285 52.295 44.300 ;
        RECT 57.300 44.285 57.630 44.300 ;
        RECT 62.625 44.285 62.955 44.300 ;
        RECT 67.960 44.285 68.290 44.300 ;
        RECT 73.285 44.285 73.615 44.300 ;
        RECT 78.620 44.285 78.950 44.300 ;
        RECT 83.945 44.285 84.275 44.300 ;
        RECT 89.280 44.285 89.610 44.300 ;
        RECT 94.605 44.285 94.935 44.300 ;
        RECT 99.940 44.285 100.270 44.300 ;
        RECT 105.265 44.285 105.595 44.300 ;
        RECT 110.600 44.285 110.930 44.300 ;
        RECT 115.925 44.285 116.255 44.300 ;
        RECT 121.260 44.285 121.590 44.300 ;
        RECT 126.585 44.285 126.915 44.300 ;
        RECT 29.705 43.985 127.180 44.285 ;
        RECT 29.735 43.970 30.935 43.985 ;
        RECT 35.980 43.970 36.310 43.985 ;
        RECT 41.305 43.970 41.635 43.985 ;
        RECT 46.640 43.970 46.970 43.985 ;
        RECT 51.965 43.970 52.295 43.985 ;
        RECT 57.300 43.970 57.630 43.985 ;
        RECT 62.625 43.970 62.955 43.985 ;
        RECT 67.960 43.970 68.290 43.985 ;
        RECT 73.285 43.970 73.615 43.985 ;
        RECT 78.620 43.970 78.950 43.985 ;
        RECT 83.945 43.970 84.275 43.985 ;
        RECT 89.280 43.970 89.610 43.985 ;
        RECT 94.605 43.970 94.935 43.985 ;
        RECT 99.940 43.970 100.270 43.985 ;
        RECT 105.265 43.970 105.595 43.985 ;
        RECT 110.600 43.970 110.930 43.985 ;
        RECT 115.925 43.970 116.255 43.985 ;
        RECT 121.260 43.970 121.590 43.985 ;
        RECT 126.585 43.970 126.915 43.985 ;
        RECT 29.735 42.950 30.935 42.965 ;
        RECT 31.480 42.950 31.810 42.965 ;
        RECT 36.805 42.950 37.135 42.965 ;
        RECT 42.140 42.950 42.470 42.965 ;
        RECT 47.465 42.950 47.795 42.965 ;
        RECT 52.800 42.950 53.130 42.965 ;
        RECT 58.125 42.950 58.455 42.965 ;
        RECT 63.460 42.950 63.790 42.965 ;
        RECT 68.785 42.950 69.115 42.965 ;
        RECT 74.120 42.950 74.450 42.965 ;
        RECT 79.445 42.950 79.775 42.965 ;
        RECT 84.780 42.950 85.110 42.965 ;
        RECT 90.105 42.950 90.435 42.965 ;
        RECT 95.440 42.950 95.770 42.965 ;
        RECT 100.765 42.950 101.095 42.965 ;
        RECT 106.100 42.950 106.430 42.965 ;
        RECT 111.425 42.950 111.755 42.965 ;
        RECT 116.760 42.950 117.090 42.965 ;
        RECT 122.085 42.950 122.415 42.965 ;
        RECT 29.705 42.650 127.180 42.950 ;
        RECT 29.735 42.635 30.935 42.650 ;
        RECT 31.480 42.635 31.810 42.650 ;
        RECT 36.805 42.635 37.135 42.650 ;
        RECT 42.140 42.635 42.470 42.650 ;
        RECT 47.465 42.635 47.795 42.650 ;
        RECT 52.800 42.635 53.130 42.650 ;
        RECT 58.125 42.635 58.455 42.650 ;
        RECT 63.460 42.635 63.790 42.650 ;
        RECT 68.785 42.635 69.115 42.650 ;
        RECT 74.120 42.635 74.450 42.650 ;
        RECT 79.445 42.635 79.775 42.650 ;
        RECT 84.780 42.635 85.110 42.650 ;
        RECT 90.105 42.635 90.435 42.650 ;
        RECT 95.440 42.635 95.770 42.650 ;
        RECT 100.765 42.635 101.095 42.650 ;
        RECT 106.100 42.635 106.430 42.650 ;
        RECT 111.425 42.635 111.755 42.650 ;
        RECT 116.760 42.635 117.090 42.650 ;
        RECT 122.085 42.635 122.415 42.650 ;
        RECT 29.735 42.305 30.935 42.320 ;
        RECT 35.980 42.305 36.310 42.320 ;
        RECT 41.305 42.305 41.635 42.320 ;
        RECT 46.640 42.305 46.970 42.320 ;
        RECT 51.965 42.305 52.295 42.320 ;
        RECT 57.300 42.305 57.630 42.320 ;
        RECT 62.625 42.305 62.955 42.320 ;
        RECT 67.960 42.305 68.290 42.320 ;
        RECT 73.285 42.305 73.615 42.320 ;
        RECT 78.620 42.305 78.950 42.320 ;
        RECT 83.945 42.305 84.275 42.320 ;
        RECT 89.280 42.305 89.610 42.320 ;
        RECT 94.605 42.305 94.935 42.320 ;
        RECT 99.940 42.305 100.270 42.320 ;
        RECT 105.265 42.305 105.595 42.320 ;
        RECT 110.600 42.305 110.930 42.320 ;
        RECT 115.925 42.305 116.255 42.320 ;
        RECT 121.260 42.305 121.590 42.320 ;
        RECT 126.585 42.305 126.915 42.320 ;
        RECT 29.705 42.005 127.180 42.305 ;
        RECT 29.735 41.990 30.935 42.005 ;
        RECT 35.980 41.990 36.310 42.005 ;
        RECT 41.305 41.990 41.635 42.005 ;
        RECT 46.640 41.990 46.970 42.005 ;
        RECT 51.965 41.990 52.295 42.005 ;
        RECT 57.300 41.990 57.630 42.005 ;
        RECT 62.625 41.990 62.955 42.005 ;
        RECT 67.960 41.990 68.290 42.005 ;
        RECT 73.285 41.990 73.615 42.005 ;
        RECT 78.620 41.990 78.950 42.005 ;
        RECT 83.945 41.990 84.275 42.005 ;
        RECT 89.280 41.990 89.610 42.005 ;
        RECT 94.605 41.990 94.935 42.005 ;
        RECT 99.940 41.990 100.270 42.005 ;
        RECT 105.265 41.990 105.595 42.005 ;
        RECT 110.600 41.990 110.930 42.005 ;
        RECT 115.925 41.990 116.255 42.005 ;
        RECT 121.260 41.990 121.590 42.005 ;
        RECT 126.585 41.990 126.915 42.005 ;
        RECT 29.735 41.660 30.935 41.675 ;
        RECT 31.480 41.660 31.810 41.670 ;
        RECT 36.805 41.660 37.135 41.670 ;
        RECT 42.140 41.660 42.470 41.670 ;
        RECT 47.465 41.660 47.795 41.670 ;
        RECT 52.800 41.660 53.130 41.670 ;
        RECT 58.125 41.660 58.455 41.670 ;
        RECT 63.460 41.660 63.790 41.670 ;
        RECT 68.785 41.660 69.115 41.670 ;
        RECT 74.120 41.660 74.450 41.670 ;
        RECT 79.445 41.660 79.775 41.670 ;
        RECT 84.780 41.660 85.110 41.670 ;
        RECT 90.105 41.660 90.435 41.670 ;
        RECT 95.440 41.660 95.770 41.670 ;
        RECT 100.765 41.660 101.095 41.670 ;
        RECT 106.100 41.660 106.430 41.670 ;
        RECT 111.425 41.660 111.755 41.670 ;
        RECT 116.760 41.660 117.090 41.670 ;
        RECT 122.085 41.660 122.415 41.670 ;
        RECT 29.705 41.360 127.180 41.660 ;
        RECT 29.735 41.345 30.935 41.360 ;
        RECT 31.480 41.340 31.810 41.360 ;
        RECT 36.805 41.340 37.135 41.360 ;
        RECT 42.140 41.340 42.470 41.360 ;
        RECT 47.465 41.340 47.795 41.360 ;
        RECT 52.800 41.340 53.130 41.360 ;
        RECT 58.125 41.340 58.455 41.360 ;
        RECT 63.460 41.340 63.790 41.360 ;
        RECT 68.785 41.340 69.115 41.360 ;
        RECT 74.120 41.340 74.450 41.360 ;
        RECT 79.445 41.340 79.775 41.360 ;
        RECT 84.780 41.340 85.110 41.360 ;
        RECT 90.105 41.340 90.435 41.360 ;
        RECT 95.440 41.340 95.770 41.360 ;
        RECT 100.765 41.340 101.095 41.360 ;
        RECT 106.100 41.340 106.430 41.360 ;
        RECT 111.425 41.340 111.755 41.360 ;
        RECT 116.760 41.340 117.090 41.360 ;
        RECT 122.085 41.340 122.415 41.360 ;
        RECT 29.735 41.015 30.935 41.030 ;
        RECT 35.985 41.015 36.315 41.040 ;
        RECT 41.310 41.015 41.640 41.040 ;
        RECT 46.645 41.015 46.975 41.040 ;
        RECT 51.970 41.015 52.300 41.040 ;
        RECT 57.305 41.015 57.635 41.040 ;
        RECT 62.630 41.015 62.960 41.040 ;
        RECT 67.965 41.015 68.295 41.040 ;
        RECT 73.290 41.015 73.620 41.040 ;
        RECT 78.625 41.015 78.955 41.040 ;
        RECT 83.950 41.015 84.280 41.040 ;
        RECT 89.285 41.015 89.615 41.040 ;
        RECT 94.610 41.015 94.940 41.040 ;
        RECT 99.945 41.015 100.275 41.040 ;
        RECT 105.270 41.015 105.600 41.040 ;
        RECT 110.605 41.015 110.935 41.040 ;
        RECT 115.930 41.015 116.260 41.040 ;
        RECT 121.265 41.015 121.595 41.040 ;
        RECT 126.590 41.015 126.920 41.040 ;
        RECT 29.705 40.715 127.180 41.015 ;
        RECT 29.735 40.700 30.935 40.715 ;
        RECT 35.985 40.710 36.315 40.715 ;
        RECT 41.310 40.710 41.640 40.715 ;
        RECT 46.645 40.710 46.975 40.715 ;
        RECT 51.970 40.710 52.300 40.715 ;
        RECT 57.305 40.710 57.635 40.715 ;
        RECT 62.630 40.710 62.960 40.715 ;
        RECT 67.965 40.710 68.295 40.715 ;
        RECT 73.290 40.710 73.620 40.715 ;
        RECT 78.625 40.710 78.955 40.715 ;
        RECT 83.950 40.710 84.280 40.715 ;
        RECT 89.285 40.710 89.615 40.715 ;
        RECT 94.610 40.710 94.940 40.715 ;
        RECT 99.945 40.710 100.275 40.715 ;
        RECT 105.270 40.710 105.600 40.715 ;
        RECT 110.605 40.710 110.935 40.715 ;
        RECT 115.930 40.710 116.260 40.715 ;
        RECT 121.265 40.710 121.595 40.715 ;
        RECT 126.590 40.710 126.920 40.715 ;
        RECT 29.735 38.685 30.935 38.700 ;
        RECT 31.485 38.685 31.815 38.700 ;
        RECT 36.810 38.685 37.140 38.700 ;
        RECT 42.145 38.685 42.475 38.700 ;
        RECT 47.470 38.685 47.800 38.700 ;
        RECT 52.805 38.685 53.135 38.700 ;
        RECT 58.130 38.685 58.460 38.700 ;
        RECT 63.465 38.685 63.795 38.700 ;
        RECT 68.790 38.685 69.120 38.700 ;
        RECT 74.125 38.685 74.455 38.700 ;
        RECT 79.450 38.685 79.780 38.700 ;
        RECT 84.785 38.685 85.115 38.700 ;
        RECT 90.110 38.685 90.440 38.700 ;
        RECT 95.445 38.685 95.775 38.700 ;
        RECT 100.770 38.685 101.100 38.700 ;
        RECT 106.105 38.685 106.435 38.700 ;
        RECT 111.430 38.685 111.760 38.700 ;
        RECT 116.765 38.685 117.095 38.700 ;
        RECT 122.090 38.685 122.420 38.700 ;
        RECT 29.705 38.385 127.180 38.685 ;
        RECT 29.735 38.370 30.935 38.385 ;
        RECT 31.485 38.370 31.815 38.385 ;
        RECT 36.810 38.370 37.140 38.385 ;
        RECT 42.145 38.370 42.475 38.385 ;
        RECT 47.470 38.370 47.800 38.385 ;
        RECT 52.805 38.370 53.135 38.385 ;
        RECT 58.130 38.370 58.460 38.385 ;
        RECT 63.465 38.370 63.795 38.385 ;
        RECT 68.790 38.370 69.120 38.385 ;
        RECT 74.125 38.370 74.455 38.385 ;
        RECT 79.450 38.370 79.780 38.385 ;
        RECT 84.785 38.370 85.115 38.385 ;
        RECT 90.110 38.370 90.440 38.385 ;
        RECT 95.445 38.370 95.775 38.385 ;
        RECT 100.770 38.370 101.100 38.385 ;
        RECT 106.105 38.370 106.435 38.385 ;
        RECT 111.430 38.370 111.760 38.385 ;
        RECT 116.765 38.370 117.095 38.385 ;
        RECT 122.090 38.370 122.420 38.385 ;
        RECT 29.735 38.040 30.935 38.055 ;
        RECT 35.980 38.040 36.310 38.055 ;
        RECT 41.305 38.040 41.635 38.055 ;
        RECT 46.640 38.040 46.970 38.055 ;
        RECT 51.965 38.040 52.295 38.055 ;
        RECT 57.300 38.040 57.630 38.055 ;
        RECT 62.625 38.040 62.955 38.055 ;
        RECT 67.960 38.040 68.290 38.055 ;
        RECT 73.285 38.040 73.615 38.055 ;
        RECT 78.620 38.040 78.950 38.055 ;
        RECT 83.945 38.040 84.275 38.055 ;
        RECT 89.280 38.040 89.610 38.055 ;
        RECT 94.605 38.040 94.935 38.055 ;
        RECT 99.940 38.040 100.270 38.055 ;
        RECT 105.265 38.040 105.595 38.055 ;
        RECT 110.600 38.040 110.930 38.055 ;
        RECT 115.925 38.040 116.255 38.055 ;
        RECT 121.260 38.040 121.590 38.055 ;
        RECT 126.585 38.040 126.915 38.055 ;
        RECT 29.705 37.740 127.180 38.040 ;
        RECT 29.735 37.725 30.935 37.740 ;
        RECT 35.980 37.725 36.310 37.740 ;
        RECT 41.305 37.725 41.635 37.740 ;
        RECT 46.640 37.725 46.970 37.740 ;
        RECT 51.965 37.725 52.295 37.740 ;
        RECT 57.300 37.725 57.630 37.740 ;
        RECT 62.625 37.725 62.955 37.740 ;
        RECT 67.960 37.725 68.290 37.740 ;
        RECT 73.285 37.725 73.615 37.740 ;
        RECT 78.620 37.725 78.950 37.740 ;
        RECT 83.945 37.725 84.275 37.740 ;
        RECT 89.280 37.725 89.610 37.740 ;
        RECT 94.605 37.725 94.935 37.740 ;
        RECT 99.940 37.725 100.270 37.740 ;
        RECT 105.265 37.725 105.595 37.740 ;
        RECT 110.600 37.725 110.930 37.740 ;
        RECT 115.925 37.725 116.255 37.740 ;
        RECT 121.260 37.725 121.590 37.740 ;
        RECT 126.585 37.725 126.915 37.740 ;
        RECT 29.735 37.395 30.935 37.410 ;
        RECT 31.480 37.395 31.810 37.410 ;
        RECT 36.805 37.395 37.135 37.410 ;
        RECT 42.140 37.395 42.470 37.410 ;
        RECT 47.465 37.395 47.795 37.410 ;
        RECT 52.800 37.395 53.130 37.410 ;
        RECT 58.125 37.395 58.455 37.410 ;
        RECT 63.460 37.395 63.790 37.410 ;
        RECT 68.785 37.395 69.115 37.410 ;
        RECT 74.120 37.395 74.450 37.410 ;
        RECT 79.445 37.395 79.775 37.410 ;
        RECT 84.780 37.395 85.110 37.410 ;
        RECT 90.105 37.395 90.435 37.410 ;
        RECT 95.440 37.395 95.770 37.410 ;
        RECT 100.765 37.395 101.095 37.410 ;
        RECT 106.100 37.395 106.430 37.410 ;
        RECT 111.425 37.395 111.755 37.410 ;
        RECT 116.760 37.395 117.090 37.410 ;
        RECT 122.085 37.395 122.415 37.410 ;
        RECT 29.705 37.095 127.180 37.395 ;
        RECT 29.735 37.080 30.935 37.095 ;
        RECT 31.480 37.080 31.810 37.095 ;
        RECT 36.805 37.080 37.135 37.095 ;
        RECT 42.140 37.080 42.470 37.095 ;
        RECT 47.465 37.080 47.795 37.095 ;
        RECT 52.800 37.080 53.130 37.095 ;
        RECT 58.125 37.080 58.455 37.095 ;
        RECT 63.460 37.080 63.790 37.095 ;
        RECT 68.785 37.080 69.115 37.095 ;
        RECT 74.120 37.080 74.450 37.095 ;
        RECT 79.445 37.080 79.775 37.095 ;
        RECT 84.780 37.080 85.110 37.095 ;
        RECT 90.105 37.080 90.435 37.095 ;
        RECT 95.440 37.080 95.770 37.095 ;
        RECT 100.765 37.080 101.095 37.095 ;
        RECT 106.100 37.080 106.430 37.095 ;
        RECT 111.425 37.080 111.755 37.095 ;
        RECT 116.760 37.080 117.090 37.095 ;
        RECT 122.085 37.080 122.415 37.095 ;
        RECT 29.735 36.750 30.935 36.765 ;
        RECT 35.980 36.750 36.310 36.765 ;
        RECT 41.305 36.750 41.635 36.765 ;
        RECT 46.640 36.750 46.970 36.765 ;
        RECT 51.965 36.750 52.295 36.765 ;
        RECT 57.300 36.750 57.630 36.765 ;
        RECT 62.625 36.750 62.955 36.765 ;
        RECT 67.960 36.750 68.290 36.765 ;
        RECT 73.285 36.750 73.615 36.765 ;
        RECT 78.620 36.750 78.950 36.765 ;
        RECT 83.945 36.750 84.275 36.765 ;
        RECT 89.280 36.750 89.610 36.765 ;
        RECT 94.605 36.750 94.935 36.765 ;
        RECT 99.940 36.750 100.270 36.765 ;
        RECT 105.265 36.750 105.595 36.765 ;
        RECT 110.600 36.750 110.930 36.765 ;
        RECT 115.925 36.750 116.255 36.765 ;
        RECT 121.260 36.750 121.590 36.765 ;
        RECT 126.585 36.750 126.915 36.765 ;
        RECT 29.705 36.450 127.180 36.750 ;
        RECT 29.735 36.435 30.935 36.450 ;
        RECT 35.980 36.435 36.310 36.450 ;
        RECT 41.305 36.435 41.635 36.450 ;
        RECT 46.640 36.435 46.970 36.450 ;
        RECT 51.965 36.435 52.295 36.450 ;
        RECT 57.300 36.435 57.630 36.450 ;
        RECT 62.625 36.435 62.955 36.450 ;
        RECT 67.960 36.435 68.290 36.450 ;
        RECT 73.285 36.435 73.615 36.450 ;
        RECT 78.620 36.435 78.950 36.450 ;
        RECT 83.945 36.435 84.275 36.450 ;
        RECT 89.280 36.435 89.610 36.450 ;
        RECT 94.605 36.435 94.935 36.450 ;
        RECT 99.940 36.435 100.270 36.450 ;
        RECT 105.265 36.435 105.595 36.450 ;
        RECT 110.600 36.435 110.930 36.450 ;
        RECT 115.925 36.435 116.255 36.450 ;
        RECT 121.260 36.435 121.590 36.450 ;
        RECT 126.585 36.435 126.915 36.450 ;
        RECT 29.735 35.415 30.935 35.430 ;
        RECT 31.480 35.415 31.810 35.430 ;
        RECT 36.805 35.415 37.135 35.430 ;
        RECT 42.140 35.415 42.470 35.430 ;
        RECT 47.465 35.415 47.795 35.430 ;
        RECT 52.800 35.415 53.130 35.430 ;
        RECT 58.125 35.415 58.455 35.430 ;
        RECT 63.460 35.415 63.790 35.430 ;
        RECT 68.785 35.415 69.115 35.430 ;
        RECT 74.120 35.415 74.450 35.430 ;
        RECT 79.445 35.415 79.775 35.430 ;
        RECT 84.780 35.415 85.110 35.430 ;
        RECT 90.105 35.415 90.435 35.430 ;
        RECT 95.440 35.415 95.770 35.430 ;
        RECT 100.765 35.415 101.095 35.430 ;
        RECT 106.100 35.415 106.430 35.430 ;
        RECT 111.425 35.415 111.755 35.430 ;
        RECT 116.760 35.415 117.090 35.430 ;
        RECT 122.085 35.415 122.415 35.430 ;
        RECT 29.705 35.115 127.180 35.415 ;
        RECT 29.735 35.100 30.935 35.115 ;
        RECT 31.480 35.100 31.810 35.115 ;
        RECT 36.805 35.100 37.135 35.115 ;
        RECT 42.140 35.100 42.470 35.115 ;
        RECT 47.465 35.100 47.795 35.115 ;
        RECT 52.800 35.100 53.130 35.115 ;
        RECT 58.125 35.100 58.455 35.115 ;
        RECT 63.460 35.100 63.790 35.115 ;
        RECT 68.785 35.100 69.115 35.115 ;
        RECT 74.120 35.100 74.450 35.115 ;
        RECT 79.445 35.100 79.775 35.115 ;
        RECT 84.780 35.100 85.110 35.115 ;
        RECT 90.105 35.100 90.435 35.115 ;
        RECT 95.440 35.100 95.770 35.115 ;
        RECT 100.765 35.100 101.095 35.115 ;
        RECT 106.100 35.100 106.430 35.115 ;
        RECT 111.425 35.100 111.755 35.115 ;
        RECT 116.760 35.100 117.090 35.115 ;
        RECT 122.085 35.100 122.415 35.115 ;
        RECT 29.735 34.770 30.935 34.785 ;
        RECT 35.980 34.770 36.310 34.785 ;
        RECT 41.305 34.770 41.635 34.785 ;
        RECT 46.640 34.770 46.970 34.785 ;
        RECT 51.965 34.770 52.295 34.785 ;
        RECT 57.300 34.770 57.630 34.785 ;
        RECT 62.625 34.770 62.955 34.785 ;
        RECT 67.960 34.770 68.290 34.785 ;
        RECT 73.285 34.770 73.615 34.785 ;
        RECT 78.620 34.770 78.950 34.785 ;
        RECT 83.945 34.770 84.275 34.785 ;
        RECT 89.280 34.770 89.610 34.785 ;
        RECT 94.605 34.770 94.935 34.785 ;
        RECT 99.940 34.770 100.270 34.785 ;
        RECT 105.265 34.770 105.595 34.785 ;
        RECT 110.600 34.770 110.930 34.785 ;
        RECT 115.925 34.770 116.255 34.785 ;
        RECT 121.260 34.770 121.590 34.785 ;
        RECT 126.585 34.770 126.915 34.785 ;
        RECT 29.705 34.470 127.180 34.770 ;
        RECT 29.735 34.455 30.935 34.470 ;
        RECT 35.980 34.455 36.310 34.470 ;
        RECT 41.305 34.455 41.635 34.470 ;
        RECT 46.640 34.455 46.970 34.470 ;
        RECT 51.965 34.455 52.295 34.470 ;
        RECT 57.300 34.455 57.630 34.470 ;
        RECT 62.625 34.455 62.955 34.470 ;
        RECT 67.960 34.455 68.290 34.470 ;
        RECT 73.285 34.455 73.615 34.470 ;
        RECT 78.620 34.455 78.950 34.470 ;
        RECT 83.945 34.455 84.275 34.470 ;
        RECT 89.280 34.455 89.610 34.470 ;
        RECT 94.605 34.455 94.935 34.470 ;
        RECT 99.940 34.455 100.270 34.470 ;
        RECT 105.265 34.455 105.595 34.470 ;
        RECT 110.600 34.455 110.930 34.470 ;
        RECT 115.925 34.455 116.255 34.470 ;
        RECT 121.260 34.455 121.590 34.470 ;
        RECT 126.585 34.455 126.915 34.470 ;
        RECT 29.735 34.125 30.935 34.140 ;
        RECT 31.480 34.125 31.810 34.135 ;
        RECT 36.805 34.125 37.135 34.135 ;
        RECT 42.140 34.125 42.470 34.135 ;
        RECT 47.465 34.125 47.795 34.135 ;
        RECT 52.800 34.125 53.130 34.135 ;
        RECT 58.125 34.125 58.455 34.135 ;
        RECT 63.460 34.125 63.790 34.135 ;
        RECT 68.785 34.125 69.115 34.135 ;
        RECT 74.120 34.125 74.450 34.135 ;
        RECT 79.445 34.125 79.775 34.135 ;
        RECT 84.780 34.125 85.110 34.135 ;
        RECT 90.105 34.125 90.435 34.135 ;
        RECT 95.440 34.125 95.770 34.135 ;
        RECT 100.765 34.125 101.095 34.135 ;
        RECT 106.100 34.125 106.430 34.135 ;
        RECT 111.425 34.125 111.755 34.135 ;
        RECT 116.760 34.125 117.090 34.135 ;
        RECT 122.085 34.125 122.415 34.135 ;
        RECT 29.705 33.825 127.180 34.125 ;
        RECT 29.735 33.810 30.935 33.825 ;
        RECT 31.480 33.805 31.810 33.825 ;
        RECT 36.805 33.805 37.135 33.825 ;
        RECT 42.140 33.805 42.470 33.825 ;
        RECT 47.465 33.805 47.795 33.825 ;
        RECT 52.800 33.805 53.130 33.825 ;
        RECT 58.125 33.805 58.455 33.825 ;
        RECT 63.460 33.805 63.790 33.825 ;
        RECT 68.785 33.805 69.115 33.825 ;
        RECT 74.120 33.805 74.450 33.825 ;
        RECT 79.445 33.805 79.775 33.825 ;
        RECT 84.780 33.805 85.110 33.825 ;
        RECT 90.105 33.805 90.435 33.825 ;
        RECT 95.440 33.805 95.770 33.825 ;
        RECT 100.765 33.805 101.095 33.825 ;
        RECT 106.100 33.805 106.430 33.825 ;
        RECT 111.425 33.805 111.755 33.825 ;
        RECT 116.760 33.805 117.090 33.825 ;
        RECT 122.085 33.805 122.415 33.825 ;
        RECT 29.735 33.480 30.935 33.495 ;
        RECT 35.985 33.480 36.315 33.505 ;
        RECT 41.310 33.480 41.640 33.505 ;
        RECT 46.645 33.480 46.975 33.505 ;
        RECT 51.970 33.480 52.300 33.505 ;
        RECT 57.305 33.480 57.635 33.505 ;
        RECT 62.630 33.480 62.960 33.505 ;
        RECT 67.965 33.480 68.295 33.505 ;
        RECT 73.290 33.480 73.620 33.505 ;
        RECT 78.625 33.480 78.955 33.505 ;
        RECT 83.950 33.480 84.280 33.505 ;
        RECT 89.285 33.480 89.615 33.505 ;
        RECT 94.610 33.480 94.940 33.505 ;
        RECT 99.945 33.480 100.275 33.505 ;
        RECT 105.270 33.480 105.600 33.505 ;
        RECT 110.605 33.480 110.935 33.505 ;
        RECT 115.930 33.480 116.260 33.505 ;
        RECT 121.265 33.480 121.595 33.505 ;
        RECT 126.590 33.480 126.920 33.505 ;
        RECT 29.705 33.180 127.180 33.480 ;
        RECT 29.735 33.165 30.935 33.180 ;
        RECT 35.985 33.175 36.315 33.180 ;
        RECT 41.310 33.175 41.640 33.180 ;
        RECT 46.645 33.175 46.975 33.180 ;
        RECT 51.970 33.175 52.300 33.180 ;
        RECT 57.305 33.175 57.635 33.180 ;
        RECT 62.630 33.175 62.960 33.180 ;
        RECT 67.965 33.175 68.295 33.180 ;
        RECT 73.290 33.175 73.620 33.180 ;
        RECT 78.625 33.175 78.955 33.180 ;
        RECT 83.950 33.175 84.280 33.180 ;
        RECT 89.285 33.175 89.615 33.180 ;
        RECT 94.610 33.175 94.940 33.180 ;
        RECT 99.945 33.175 100.275 33.180 ;
        RECT 105.270 33.175 105.600 33.180 ;
        RECT 110.605 33.175 110.935 33.180 ;
        RECT 115.930 33.175 116.260 33.180 ;
        RECT 121.265 33.175 121.595 33.180 ;
        RECT 126.590 33.175 126.920 33.180 ;
        RECT 29.735 31.150 30.935 31.165 ;
        RECT 31.485 31.150 31.815 31.165 ;
        RECT 36.810 31.150 37.140 31.165 ;
        RECT 42.145 31.150 42.475 31.165 ;
        RECT 47.470 31.150 47.800 31.165 ;
        RECT 52.805 31.150 53.135 31.165 ;
        RECT 58.130 31.150 58.460 31.165 ;
        RECT 63.465 31.150 63.795 31.165 ;
        RECT 68.790 31.150 69.120 31.165 ;
        RECT 74.125 31.150 74.455 31.165 ;
        RECT 79.450 31.150 79.780 31.165 ;
        RECT 84.785 31.150 85.115 31.165 ;
        RECT 90.110 31.150 90.440 31.165 ;
        RECT 95.445 31.150 95.775 31.165 ;
        RECT 100.770 31.150 101.100 31.165 ;
        RECT 106.105 31.150 106.435 31.165 ;
        RECT 111.430 31.150 111.760 31.165 ;
        RECT 116.765 31.150 117.095 31.165 ;
        RECT 122.090 31.150 122.420 31.165 ;
        RECT 29.705 30.850 127.180 31.150 ;
        RECT 29.735 30.835 30.935 30.850 ;
        RECT 31.485 30.835 31.815 30.850 ;
        RECT 36.810 30.835 37.140 30.850 ;
        RECT 42.145 30.835 42.475 30.850 ;
        RECT 47.470 30.835 47.800 30.850 ;
        RECT 52.805 30.835 53.135 30.850 ;
        RECT 58.130 30.835 58.460 30.850 ;
        RECT 63.465 30.835 63.795 30.850 ;
        RECT 68.790 30.835 69.120 30.850 ;
        RECT 74.125 30.835 74.455 30.850 ;
        RECT 79.450 30.835 79.780 30.850 ;
        RECT 84.785 30.835 85.115 30.850 ;
        RECT 90.110 30.835 90.440 30.850 ;
        RECT 95.445 30.835 95.775 30.850 ;
        RECT 100.770 30.835 101.100 30.850 ;
        RECT 106.105 30.835 106.435 30.850 ;
        RECT 111.430 30.835 111.760 30.850 ;
        RECT 116.765 30.835 117.095 30.850 ;
        RECT 122.090 30.835 122.420 30.850 ;
        RECT 29.735 30.505 30.935 30.520 ;
        RECT 35.980 30.505 36.310 30.520 ;
        RECT 41.305 30.505 41.635 30.520 ;
        RECT 46.640 30.505 46.970 30.520 ;
        RECT 51.965 30.505 52.295 30.520 ;
        RECT 57.300 30.505 57.630 30.520 ;
        RECT 62.625 30.505 62.955 30.520 ;
        RECT 67.960 30.505 68.290 30.520 ;
        RECT 73.285 30.505 73.615 30.520 ;
        RECT 78.620 30.505 78.950 30.520 ;
        RECT 83.945 30.505 84.275 30.520 ;
        RECT 89.280 30.505 89.610 30.520 ;
        RECT 94.605 30.505 94.935 30.520 ;
        RECT 99.940 30.505 100.270 30.520 ;
        RECT 105.265 30.505 105.595 30.520 ;
        RECT 110.600 30.505 110.930 30.520 ;
        RECT 115.925 30.505 116.255 30.520 ;
        RECT 121.260 30.505 121.590 30.520 ;
        RECT 126.585 30.505 126.915 30.520 ;
        RECT 29.705 30.205 127.180 30.505 ;
        RECT 29.735 30.190 30.935 30.205 ;
        RECT 35.980 30.190 36.310 30.205 ;
        RECT 41.305 30.190 41.635 30.205 ;
        RECT 46.640 30.190 46.970 30.205 ;
        RECT 51.965 30.190 52.295 30.205 ;
        RECT 57.300 30.190 57.630 30.205 ;
        RECT 62.625 30.190 62.955 30.205 ;
        RECT 67.960 30.190 68.290 30.205 ;
        RECT 73.285 30.190 73.615 30.205 ;
        RECT 78.620 30.190 78.950 30.205 ;
        RECT 83.945 30.190 84.275 30.205 ;
        RECT 89.280 30.190 89.610 30.205 ;
        RECT 94.605 30.190 94.935 30.205 ;
        RECT 99.940 30.190 100.270 30.205 ;
        RECT 105.265 30.190 105.595 30.205 ;
        RECT 110.600 30.190 110.930 30.205 ;
        RECT 115.925 30.190 116.255 30.205 ;
        RECT 121.260 30.190 121.590 30.205 ;
        RECT 126.585 30.190 126.915 30.205 ;
        RECT 29.735 29.860 30.935 29.875 ;
        RECT 31.480 29.860 31.810 29.875 ;
        RECT 36.805 29.860 37.135 29.875 ;
        RECT 42.140 29.860 42.470 29.875 ;
        RECT 47.465 29.860 47.795 29.875 ;
        RECT 52.800 29.860 53.130 29.875 ;
        RECT 58.125 29.860 58.455 29.875 ;
        RECT 63.460 29.860 63.790 29.875 ;
        RECT 68.785 29.860 69.115 29.875 ;
        RECT 74.120 29.860 74.450 29.875 ;
        RECT 79.445 29.860 79.775 29.875 ;
        RECT 84.780 29.860 85.110 29.875 ;
        RECT 90.105 29.860 90.435 29.875 ;
        RECT 95.440 29.860 95.770 29.875 ;
        RECT 100.765 29.860 101.095 29.875 ;
        RECT 106.100 29.860 106.430 29.875 ;
        RECT 111.425 29.860 111.755 29.875 ;
        RECT 116.760 29.860 117.090 29.875 ;
        RECT 122.085 29.860 122.415 29.875 ;
        RECT 29.705 29.560 127.180 29.860 ;
        RECT 29.735 29.545 30.935 29.560 ;
        RECT 31.480 29.545 31.810 29.560 ;
        RECT 36.805 29.545 37.135 29.560 ;
        RECT 42.140 29.545 42.470 29.560 ;
        RECT 47.465 29.545 47.795 29.560 ;
        RECT 52.800 29.545 53.130 29.560 ;
        RECT 58.125 29.545 58.455 29.560 ;
        RECT 63.460 29.545 63.790 29.560 ;
        RECT 68.785 29.545 69.115 29.560 ;
        RECT 74.120 29.545 74.450 29.560 ;
        RECT 79.445 29.545 79.775 29.560 ;
        RECT 84.780 29.545 85.110 29.560 ;
        RECT 90.105 29.545 90.435 29.560 ;
        RECT 95.440 29.545 95.770 29.560 ;
        RECT 100.765 29.545 101.095 29.560 ;
        RECT 106.100 29.545 106.430 29.560 ;
        RECT 111.425 29.545 111.755 29.560 ;
        RECT 116.760 29.545 117.090 29.560 ;
        RECT 122.085 29.545 122.415 29.560 ;
        RECT 29.735 29.215 30.935 29.230 ;
        RECT 35.980 29.215 36.310 29.230 ;
        RECT 41.305 29.215 41.635 29.230 ;
        RECT 46.640 29.215 46.970 29.230 ;
        RECT 51.965 29.215 52.295 29.230 ;
        RECT 57.300 29.215 57.630 29.230 ;
        RECT 62.625 29.215 62.955 29.230 ;
        RECT 67.960 29.215 68.290 29.230 ;
        RECT 73.285 29.215 73.615 29.230 ;
        RECT 78.620 29.215 78.950 29.230 ;
        RECT 83.945 29.215 84.275 29.230 ;
        RECT 89.280 29.215 89.610 29.230 ;
        RECT 94.605 29.215 94.935 29.230 ;
        RECT 99.940 29.215 100.270 29.230 ;
        RECT 105.265 29.215 105.595 29.230 ;
        RECT 110.600 29.215 110.930 29.230 ;
        RECT 115.925 29.215 116.255 29.230 ;
        RECT 121.260 29.215 121.590 29.230 ;
        RECT 126.585 29.215 126.915 29.230 ;
        RECT 29.705 28.915 127.180 29.215 ;
        RECT 29.735 28.900 30.935 28.915 ;
        RECT 35.980 28.900 36.310 28.915 ;
        RECT 41.305 28.900 41.635 28.915 ;
        RECT 46.640 28.900 46.970 28.915 ;
        RECT 51.965 28.900 52.295 28.915 ;
        RECT 57.300 28.900 57.630 28.915 ;
        RECT 62.625 28.900 62.955 28.915 ;
        RECT 67.960 28.900 68.290 28.915 ;
        RECT 73.285 28.900 73.615 28.915 ;
        RECT 78.620 28.900 78.950 28.915 ;
        RECT 83.945 28.900 84.275 28.915 ;
        RECT 89.280 28.900 89.610 28.915 ;
        RECT 94.605 28.900 94.935 28.915 ;
        RECT 99.940 28.900 100.270 28.915 ;
        RECT 105.265 28.900 105.595 28.915 ;
        RECT 110.600 28.900 110.930 28.915 ;
        RECT 115.925 28.900 116.255 28.915 ;
        RECT 121.260 28.900 121.590 28.915 ;
        RECT 126.585 28.900 126.915 28.915 ;
        RECT 29.735 27.880 30.935 27.895 ;
        RECT 31.480 27.880 31.810 27.895 ;
        RECT 36.805 27.880 37.135 27.895 ;
        RECT 42.140 27.880 42.470 27.895 ;
        RECT 47.465 27.880 47.795 27.895 ;
        RECT 52.800 27.880 53.130 27.895 ;
        RECT 58.125 27.880 58.455 27.895 ;
        RECT 63.460 27.880 63.790 27.895 ;
        RECT 68.785 27.880 69.115 27.895 ;
        RECT 74.120 27.880 74.450 27.895 ;
        RECT 79.445 27.880 79.775 27.895 ;
        RECT 84.780 27.880 85.110 27.895 ;
        RECT 90.105 27.880 90.435 27.895 ;
        RECT 95.440 27.880 95.770 27.895 ;
        RECT 100.765 27.880 101.095 27.895 ;
        RECT 106.100 27.880 106.430 27.895 ;
        RECT 111.425 27.880 111.755 27.895 ;
        RECT 116.760 27.880 117.090 27.895 ;
        RECT 122.085 27.880 122.415 27.895 ;
        RECT 29.705 27.580 127.180 27.880 ;
        RECT 29.735 27.565 30.935 27.580 ;
        RECT 31.480 27.565 31.810 27.580 ;
        RECT 36.805 27.565 37.135 27.580 ;
        RECT 42.140 27.565 42.470 27.580 ;
        RECT 47.465 27.565 47.795 27.580 ;
        RECT 52.800 27.565 53.130 27.580 ;
        RECT 58.125 27.565 58.455 27.580 ;
        RECT 63.460 27.565 63.790 27.580 ;
        RECT 68.785 27.565 69.115 27.580 ;
        RECT 74.120 27.565 74.450 27.580 ;
        RECT 79.445 27.565 79.775 27.580 ;
        RECT 84.780 27.565 85.110 27.580 ;
        RECT 90.105 27.565 90.435 27.580 ;
        RECT 95.440 27.565 95.770 27.580 ;
        RECT 100.765 27.565 101.095 27.580 ;
        RECT 106.100 27.565 106.430 27.580 ;
        RECT 111.425 27.565 111.755 27.580 ;
        RECT 116.760 27.565 117.090 27.580 ;
        RECT 122.085 27.565 122.415 27.580 ;
        RECT 29.735 27.235 30.935 27.250 ;
        RECT 35.980 27.235 36.310 27.250 ;
        RECT 41.305 27.235 41.635 27.250 ;
        RECT 46.640 27.235 46.970 27.250 ;
        RECT 51.965 27.235 52.295 27.250 ;
        RECT 57.300 27.235 57.630 27.250 ;
        RECT 62.625 27.235 62.955 27.250 ;
        RECT 67.960 27.235 68.290 27.250 ;
        RECT 73.285 27.235 73.615 27.250 ;
        RECT 78.620 27.235 78.950 27.250 ;
        RECT 83.945 27.235 84.275 27.250 ;
        RECT 89.280 27.235 89.610 27.250 ;
        RECT 94.605 27.235 94.935 27.250 ;
        RECT 99.940 27.235 100.270 27.250 ;
        RECT 105.265 27.235 105.595 27.250 ;
        RECT 110.600 27.235 110.930 27.250 ;
        RECT 115.925 27.235 116.255 27.250 ;
        RECT 121.260 27.235 121.590 27.250 ;
        RECT 126.585 27.235 126.915 27.250 ;
        RECT 29.705 26.935 127.180 27.235 ;
        RECT 29.735 26.920 30.935 26.935 ;
        RECT 35.980 26.920 36.310 26.935 ;
        RECT 41.305 26.920 41.635 26.935 ;
        RECT 46.640 26.920 46.970 26.935 ;
        RECT 51.965 26.920 52.295 26.935 ;
        RECT 57.300 26.920 57.630 26.935 ;
        RECT 62.625 26.920 62.955 26.935 ;
        RECT 67.960 26.920 68.290 26.935 ;
        RECT 73.285 26.920 73.615 26.935 ;
        RECT 78.620 26.920 78.950 26.935 ;
        RECT 83.945 26.920 84.275 26.935 ;
        RECT 89.280 26.920 89.610 26.935 ;
        RECT 94.605 26.920 94.935 26.935 ;
        RECT 99.940 26.920 100.270 26.935 ;
        RECT 105.265 26.920 105.595 26.935 ;
        RECT 110.600 26.920 110.930 26.935 ;
        RECT 115.925 26.920 116.255 26.935 ;
        RECT 121.260 26.920 121.590 26.935 ;
        RECT 126.585 26.920 126.915 26.935 ;
        RECT 29.735 26.590 30.935 26.605 ;
        RECT 31.480 26.590 31.810 26.600 ;
        RECT 36.805 26.590 37.135 26.600 ;
        RECT 42.140 26.590 42.470 26.600 ;
        RECT 47.465 26.590 47.795 26.600 ;
        RECT 52.800 26.590 53.130 26.600 ;
        RECT 58.125 26.590 58.455 26.600 ;
        RECT 63.460 26.590 63.790 26.600 ;
        RECT 68.785 26.590 69.115 26.600 ;
        RECT 74.120 26.590 74.450 26.600 ;
        RECT 79.445 26.590 79.775 26.600 ;
        RECT 84.780 26.590 85.110 26.600 ;
        RECT 90.105 26.590 90.435 26.600 ;
        RECT 95.440 26.590 95.770 26.600 ;
        RECT 100.765 26.590 101.095 26.600 ;
        RECT 106.100 26.590 106.430 26.600 ;
        RECT 111.425 26.590 111.755 26.600 ;
        RECT 116.760 26.590 117.090 26.600 ;
        RECT 122.085 26.590 122.415 26.600 ;
        RECT 29.705 26.290 127.180 26.590 ;
        RECT 29.735 26.275 30.935 26.290 ;
        RECT 31.480 26.270 31.810 26.290 ;
        RECT 36.805 26.270 37.135 26.290 ;
        RECT 42.140 26.270 42.470 26.290 ;
        RECT 47.465 26.270 47.795 26.290 ;
        RECT 52.800 26.270 53.130 26.290 ;
        RECT 58.125 26.270 58.455 26.290 ;
        RECT 63.460 26.270 63.790 26.290 ;
        RECT 68.785 26.270 69.115 26.290 ;
        RECT 74.120 26.270 74.450 26.290 ;
        RECT 79.445 26.270 79.775 26.290 ;
        RECT 84.780 26.270 85.110 26.290 ;
        RECT 90.105 26.270 90.435 26.290 ;
        RECT 95.440 26.270 95.770 26.290 ;
        RECT 100.765 26.270 101.095 26.290 ;
        RECT 106.100 26.270 106.430 26.290 ;
        RECT 111.425 26.270 111.755 26.290 ;
        RECT 116.760 26.270 117.090 26.290 ;
        RECT 122.085 26.270 122.415 26.290 ;
        RECT 29.735 25.945 30.935 25.960 ;
        RECT 35.985 25.945 36.315 25.970 ;
        RECT 41.310 25.945 41.640 25.970 ;
        RECT 46.645 25.945 46.975 25.970 ;
        RECT 51.970 25.945 52.300 25.970 ;
        RECT 57.305 25.945 57.635 25.970 ;
        RECT 62.630 25.945 62.960 25.970 ;
        RECT 67.965 25.945 68.295 25.970 ;
        RECT 73.290 25.945 73.620 25.970 ;
        RECT 78.625 25.945 78.955 25.970 ;
        RECT 83.950 25.945 84.280 25.970 ;
        RECT 89.285 25.945 89.615 25.970 ;
        RECT 94.610 25.945 94.940 25.970 ;
        RECT 99.945 25.945 100.275 25.970 ;
        RECT 105.270 25.945 105.600 25.970 ;
        RECT 110.605 25.945 110.935 25.970 ;
        RECT 115.930 25.945 116.260 25.970 ;
        RECT 121.265 25.945 121.595 25.970 ;
        RECT 126.590 25.945 126.920 25.970 ;
        RECT 29.705 25.645 127.180 25.945 ;
        RECT 29.735 25.630 30.935 25.645 ;
        RECT 35.985 25.640 36.315 25.645 ;
        RECT 41.310 25.640 41.640 25.645 ;
        RECT 46.645 25.640 46.975 25.645 ;
        RECT 51.970 25.640 52.300 25.645 ;
        RECT 57.305 25.640 57.635 25.645 ;
        RECT 62.630 25.640 62.960 25.645 ;
        RECT 67.965 25.640 68.295 25.645 ;
        RECT 73.290 25.640 73.620 25.645 ;
        RECT 78.625 25.640 78.955 25.645 ;
        RECT 83.950 25.640 84.280 25.645 ;
        RECT 89.285 25.640 89.615 25.645 ;
        RECT 94.610 25.640 94.940 25.645 ;
        RECT 99.945 25.640 100.275 25.645 ;
        RECT 105.270 25.640 105.600 25.645 ;
        RECT 110.605 25.640 110.935 25.645 ;
        RECT 115.930 25.640 116.260 25.645 ;
        RECT 121.265 25.640 121.595 25.645 ;
        RECT 126.590 25.640 126.920 25.645 ;
        RECT 29.735 23.615 30.935 23.630 ;
        RECT 31.485 23.615 31.815 23.630 ;
        RECT 36.810 23.615 37.140 23.630 ;
        RECT 42.145 23.615 42.475 23.630 ;
        RECT 47.470 23.615 47.800 23.630 ;
        RECT 52.805 23.615 53.135 23.630 ;
        RECT 58.130 23.615 58.460 23.630 ;
        RECT 63.465 23.615 63.795 23.630 ;
        RECT 68.790 23.615 69.120 23.630 ;
        RECT 74.125 23.615 74.455 23.630 ;
        RECT 79.450 23.615 79.780 23.630 ;
        RECT 84.785 23.615 85.115 23.630 ;
        RECT 90.110 23.615 90.440 23.630 ;
        RECT 95.445 23.615 95.775 23.630 ;
        RECT 100.770 23.615 101.100 23.630 ;
        RECT 106.105 23.615 106.435 23.630 ;
        RECT 111.430 23.615 111.760 23.630 ;
        RECT 116.765 23.615 117.095 23.630 ;
        RECT 122.090 23.615 122.420 23.630 ;
        RECT 29.705 23.315 127.180 23.615 ;
        RECT 29.735 23.300 30.935 23.315 ;
        RECT 31.485 23.300 31.815 23.315 ;
        RECT 36.810 23.300 37.140 23.315 ;
        RECT 42.145 23.300 42.475 23.315 ;
        RECT 47.470 23.300 47.800 23.315 ;
        RECT 52.805 23.300 53.135 23.315 ;
        RECT 58.130 23.300 58.460 23.315 ;
        RECT 63.465 23.300 63.795 23.315 ;
        RECT 68.790 23.300 69.120 23.315 ;
        RECT 74.125 23.300 74.455 23.315 ;
        RECT 79.450 23.300 79.780 23.315 ;
        RECT 84.785 23.300 85.115 23.315 ;
        RECT 90.110 23.300 90.440 23.315 ;
        RECT 95.445 23.300 95.775 23.315 ;
        RECT 100.770 23.300 101.100 23.315 ;
        RECT 106.105 23.300 106.435 23.315 ;
        RECT 111.430 23.300 111.760 23.315 ;
        RECT 116.765 23.300 117.095 23.315 ;
        RECT 122.090 23.300 122.420 23.315 ;
        RECT 29.735 22.970 30.935 22.985 ;
        RECT 35.980 22.970 36.310 22.985 ;
        RECT 41.305 22.970 41.635 22.985 ;
        RECT 46.640 22.970 46.970 22.985 ;
        RECT 51.965 22.970 52.295 22.985 ;
        RECT 57.300 22.970 57.630 22.985 ;
        RECT 62.625 22.970 62.955 22.985 ;
        RECT 67.960 22.970 68.290 22.985 ;
        RECT 73.285 22.970 73.615 22.985 ;
        RECT 78.620 22.970 78.950 22.985 ;
        RECT 83.945 22.970 84.275 22.985 ;
        RECT 89.280 22.970 89.610 22.985 ;
        RECT 94.605 22.970 94.935 22.985 ;
        RECT 99.940 22.970 100.270 22.985 ;
        RECT 105.265 22.970 105.595 22.985 ;
        RECT 110.600 22.970 110.930 22.985 ;
        RECT 115.925 22.970 116.255 22.985 ;
        RECT 121.260 22.970 121.590 22.985 ;
        RECT 126.585 22.970 126.915 22.985 ;
        RECT 29.705 22.670 127.180 22.970 ;
        RECT 29.735 22.655 30.935 22.670 ;
        RECT 35.980 22.655 36.310 22.670 ;
        RECT 41.305 22.655 41.635 22.670 ;
        RECT 46.640 22.655 46.970 22.670 ;
        RECT 51.965 22.655 52.295 22.670 ;
        RECT 57.300 22.655 57.630 22.670 ;
        RECT 62.625 22.655 62.955 22.670 ;
        RECT 67.960 22.655 68.290 22.670 ;
        RECT 73.285 22.655 73.615 22.670 ;
        RECT 78.620 22.655 78.950 22.670 ;
        RECT 83.945 22.655 84.275 22.670 ;
        RECT 89.280 22.655 89.610 22.670 ;
        RECT 94.605 22.655 94.935 22.670 ;
        RECT 99.940 22.655 100.270 22.670 ;
        RECT 105.265 22.655 105.595 22.670 ;
        RECT 110.600 22.655 110.930 22.670 ;
        RECT 115.925 22.655 116.255 22.670 ;
        RECT 121.260 22.655 121.590 22.670 ;
        RECT 126.585 22.655 126.915 22.670 ;
        RECT 29.735 22.325 30.935 22.340 ;
        RECT 31.480 22.325 31.810 22.340 ;
        RECT 36.805 22.325 37.135 22.340 ;
        RECT 42.140 22.325 42.470 22.340 ;
        RECT 47.465 22.325 47.795 22.340 ;
        RECT 52.800 22.325 53.130 22.340 ;
        RECT 58.125 22.325 58.455 22.340 ;
        RECT 63.460 22.325 63.790 22.340 ;
        RECT 68.785 22.325 69.115 22.340 ;
        RECT 74.120 22.325 74.450 22.340 ;
        RECT 79.445 22.325 79.775 22.340 ;
        RECT 84.780 22.325 85.110 22.340 ;
        RECT 90.105 22.325 90.435 22.340 ;
        RECT 95.440 22.325 95.770 22.340 ;
        RECT 100.765 22.325 101.095 22.340 ;
        RECT 106.100 22.325 106.430 22.340 ;
        RECT 111.425 22.325 111.755 22.340 ;
        RECT 116.760 22.325 117.090 22.340 ;
        RECT 122.085 22.325 122.415 22.340 ;
        RECT 29.705 22.025 127.180 22.325 ;
        RECT 29.735 22.010 30.935 22.025 ;
        RECT 31.480 22.010 31.810 22.025 ;
        RECT 36.805 22.010 37.135 22.025 ;
        RECT 42.140 22.010 42.470 22.025 ;
        RECT 47.465 22.010 47.795 22.025 ;
        RECT 52.800 22.010 53.130 22.025 ;
        RECT 58.125 22.010 58.455 22.025 ;
        RECT 63.460 22.010 63.790 22.025 ;
        RECT 68.785 22.010 69.115 22.025 ;
        RECT 74.120 22.010 74.450 22.025 ;
        RECT 79.445 22.010 79.775 22.025 ;
        RECT 84.780 22.010 85.110 22.025 ;
        RECT 90.105 22.010 90.435 22.025 ;
        RECT 95.440 22.010 95.770 22.025 ;
        RECT 100.765 22.010 101.095 22.025 ;
        RECT 106.100 22.010 106.430 22.025 ;
        RECT 111.425 22.010 111.755 22.025 ;
        RECT 116.760 22.010 117.090 22.025 ;
        RECT 122.085 22.010 122.415 22.025 ;
        RECT 29.735 21.680 30.935 21.695 ;
        RECT 35.980 21.680 36.310 21.695 ;
        RECT 41.305 21.680 41.635 21.695 ;
        RECT 46.640 21.680 46.970 21.695 ;
        RECT 51.965 21.680 52.295 21.695 ;
        RECT 57.300 21.680 57.630 21.695 ;
        RECT 62.625 21.680 62.955 21.695 ;
        RECT 67.960 21.680 68.290 21.695 ;
        RECT 73.285 21.680 73.615 21.695 ;
        RECT 78.620 21.680 78.950 21.695 ;
        RECT 83.945 21.680 84.275 21.695 ;
        RECT 89.280 21.680 89.610 21.695 ;
        RECT 94.605 21.680 94.935 21.695 ;
        RECT 99.940 21.680 100.270 21.695 ;
        RECT 105.265 21.680 105.595 21.695 ;
        RECT 110.600 21.680 110.930 21.695 ;
        RECT 115.925 21.680 116.255 21.695 ;
        RECT 121.260 21.680 121.590 21.695 ;
        RECT 126.585 21.680 126.915 21.695 ;
        RECT 29.705 21.380 127.180 21.680 ;
        RECT 29.735 21.365 30.935 21.380 ;
        RECT 35.980 21.365 36.310 21.380 ;
        RECT 41.305 21.365 41.635 21.380 ;
        RECT 46.640 21.365 46.970 21.380 ;
        RECT 51.965 21.365 52.295 21.380 ;
        RECT 57.300 21.365 57.630 21.380 ;
        RECT 62.625 21.365 62.955 21.380 ;
        RECT 67.960 21.365 68.290 21.380 ;
        RECT 73.285 21.365 73.615 21.380 ;
        RECT 78.620 21.365 78.950 21.380 ;
        RECT 83.945 21.365 84.275 21.380 ;
        RECT 89.280 21.365 89.610 21.380 ;
        RECT 94.605 21.365 94.935 21.380 ;
        RECT 99.940 21.365 100.270 21.380 ;
        RECT 105.265 21.365 105.595 21.380 ;
        RECT 110.600 21.365 110.930 21.380 ;
        RECT 115.925 21.365 116.255 21.380 ;
        RECT 121.260 21.365 121.590 21.380 ;
        RECT 126.585 21.365 126.915 21.380 ;
        RECT 29.735 20.345 30.935 20.360 ;
        RECT 31.480 20.345 31.810 20.360 ;
        RECT 36.805 20.345 37.135 20.360 ;
        RECT 42.140 20.345 42.470 20.360 ;
        RECT 47.465 20.345 47.795 20.360 ;
        RECT 52.800 20.345 53.130 20.360 ;
        RECT 58.125 20.345 58.455 20.360 ;
        RECT 63.460 20.345 63.790 20.360 ;
        RECT 68.785 20.345 69.115 20.360 ;
        RECT 74.120 20.345 74.450 20.360 ;
        RECT 79.445 20.345 79.775 20.360 ;
        RECT 84.780 20.345 85.110 20.360 ;
        RECT 90.105 20.345 90.435 20.360 ;
        RECT 95.440 20.345 95.770 20.360 ;
        RECT 100.765 20.345 101.095 20.360 ;
        RECT 106.100 20.345 106.430 20.360 ;
        RECT 111.425 20.345 111.755 20.360 ;
        RECT 116.760 20.345 117.090 20.360 ;
        RECT 122.085 20.345 122.415 20.360 ;
        RECT 29.705 20.045 127.180 20.345 ;
        RECT 29.735 20.030 30.935 20.045 ;
        RECT 31.480 20.030 31.810 20.045 ;
        RECT 36.805 20.030 37.135 20.045 ;
        RECT 42.140 20.030 42.470 20.045 ;
        RECT 47.465 20.030 47.795 20.045 ;
        RECT 52.800 20.030 53.130 20.045 ;
        RECT 58.125 20.030 58.455 20.045 ;
        RECT 63.460 20.030 63.790 20.045 ;
        RECT 68.785 20.030 69.115 20.045 ;
        RECT 74.120 20.030 74.450 20.045 ;
        RECT 79.445 20.030 79.775 20.045 ;
        RECT 84.780 20.030 85.110 20.045 ;
        RECT 90.105 20.030 90.435 20.045 ;
        RECT 95.440 20.030 95.770 20.045 ;
        RECT 100.765 20.030 101.095 20.045 ;
        RECT 106.100 20.030 106.430 20.045 ;
        RECT 111.425 20.030 111.755 20.045 ;
        RECT 116.760 20.030 117.090 20.045 ;
        RECT 122.085 20.030 122.415 20.045 ;
        RECT 29.735 19.700 30.935 19.715 ;
        RECT 35.980 19.700 36.310 19.715 ;
        RECT 41.305 19.700 41.635 19.715 ;
        RECT 46.640 19.700 46.970 19.715 ;
        RECT 51.965 19.700 52.295 19.715 ;
        RECT 57.300 19.700 57.630 19.715 ;
        RECT 62.625 19.700 62.955 19.715 ;
        RECT 67.960 19.700 68.290 19.715 ;
        RECT 73.285 19.700 73.615 19.715 ;
        RECT 78.620 19.700 78.950 19.715 ;
        RECT 83.945 19.700 84.275 19.715 ;
        RECT 89.280 19.700 89.610 19.715 ;
        RECT 94.605 19.700 94.935 19.715 ;
        RECT 99.940 19.700 100.270 19.715 ;
        RECT 105.265 19.700 105.595 19.715 ;
        RECT 110.600 19.700 110.930 19.715 ;
        RECT 115.925 19.700 116.255 19.715 ;
        RECT 121.260 19.700 121.590 19.715 ;
        RECT 126.585 19.700 126.915 19.715 ;
        RECT 29.705 19.400 127.180 19.700 ;
        RECT 29.735 19.385 30.935 19.400 ;
        RECT 35.980 19.385 36.310 19.400 ;
        RECT 41.305 19.385 41.635 19.400 ;
        RECT 46.640 19.385 46.970 19.400 ;
        RECT 51.965 19.385 52.295 19.400 ;
        RECT 57.300 19.385 57.630 19.400 ;
        RECT 62.625 19.385 62.955 19.400 ;
        RECT 67.960 19.385 68.290 19.400 ;
        RECT 73.285 19.385 73.615 19.400 ;
        RECT 78.620 19.385 78.950 19.400 ;
        RECT 83.945 19.385 84.275 19.400 ;
        RECT 89.280 19.385 89.610 19.400 ;
        RECT 94.605 19.385 94.935 19.400 ;
        RECT 99.940 19.385 100.270 19.400 ;
        RECT 105.265 19.385 105.595 19.400 ;
        RECT 110.600 19.385 110.930 19.400 ;
        RECT 115.925 19.385 116.255 19.400 ;
        RECT 121.260 19.385 121.590 19.400 ;
        RECT 126.585 19.385 126.915 19.400 ;
        RECT 29.735 19.055 30.935 19.070 ;
        RECT 31.480 19.055 31.810 19.065 ;
        RECT 36.805 19.055 37.135 19.065 ;
        RECT 42.140 19.055 42.470 19.065 ;
        RECT 47.465 19.055 47.795 19.065 ;
        RECT 52.800 19.055 53.130 19.065 ;
        RECT 58.125 19.055 58.455 19.065 ;
        RECT 63.460 19.055 63.790 19.065 ;
        RECT 68.785 19.055 69.115 19.065 ;
        RECT 74.120 19.055 74.450 19.065 ;
        RECT 79.445 19.055 79.775 19.065 ;
        RECT 84.780 19.055 85.110 19.065 ;
        RECT 90.105 19.055 90.435 19.065 ;
        RECT 95.440 19.055 95.770 19.065 ;
        RECT 100.765 19.055 101.095 19.065 ;
        RECT 106.100 19.055 106.430 19.065 ;
        RECT 111.425 19.055 111.755 19.065 ;
        RECT 116.760 19.055 117.090 19.065 ;
        RECT 122.085 19.055 122.415 19.065 ;
        RECT 29.705 18.755 127.180 19.055 ;
        RECT 29.735 18.740 30.935 18.755 ;
        RECT 31.480 18.735 31.810 18.755 ;
        RECT 36.805 18.735 37.135 18.755 ;
        RECT 42.140 18.735 42.470 18.755 ;
        RECT 47.465 18.735 47.795 18.755 ;
        RECT 52.800 18.735 53.130 18.755 ;
        RECT 58.125 18.735 58.455 18.755 ;
        RECT 63.460 18.735 63.790 18.755 ;
        RECT 68.785 18.735 69.115 18.755 ;
        RECT 74.120 18.735 74.450 18.755 ;
        RECT 79.445 18.735 79.775 18.755 ;
        RECT 84.780 18.735 85.110 18.755 ;
        RECT 90.105 18.735 90.435 18.755 ;
        RECT 95.440 18.735 95.770 18.755 ;
        RECT 100.765 18.735 101.095 18.755 ;
        RECT 106.100 18.735 106.430 18.755 ;
        RECT 111.425 18.735 111.755 18.755 ;
        RECT 116.760 18.735 117.090 18.755 ;
        RECT 122.085 18.735 122.415 18.755 ;
        RECT 29.735 18.410 30.935 18.425 ;
        RECT 35.985 18.410 36.315 18.435 ;
        RECT 41.310 18.410 41.640 18.435 ;
        RECT 46.645 18.410 46.975 18.435 ;
        RECT 51.970 18.410 52.300 18.435 ;
        RECT 57.305 18.410 57.635 18.435 ;
        RECT 62.630 18.410 62.960 18.435 ;
        RECT 67.965 18.410 68.295 18.435 ;
        RECT 73.290 18.410 73.620 18.435 ;
        RECT 78.625 18.410 78.955 18.435 ;
        RECT 83.950 18.410 84.280 18.435 ;
        RECT 89.285 18.410 89.615 18.435 ;
        RECT 94.610 18.410 94.940 18.435 ;
        RECT 99.945 18.410 100.275 18.435 ;
        RECT 105.270 18.410 105.600 18.435 ;
        RECT 110.605 18.410 110.935 18.435 ;
        RECT 115.930 18.410 116.260 18.435 ;
        RECT 121.265 18.410 121.595 18.435 ;
        RECT 126.590 18.410 126.920 18.435 ;
        RECT 29.705 18.110 127.180 18.410 ;
        RECT 29.735 18.095 30.935 18.110 ;
        RECT 35.985 18.105 36.315 18.110 ;
        RECT 41.310 18.105 41.640 18.110 ;
        RECT 46.645 18.105 46.975 18.110 ;
        RECT 51.970 18.105 52.300 18.110 ;
        RECT 57.305 18.105 57.635 18.110 ;
        RECT 62.630 18.105 62.960 18.110 ;
        RECT 67.965 18.105 68.295 18.110 ;
        RECT 73.290 18.105 73.620 18.110 ;
        RECT 78.625 18.105 78.955 18.110 ;
        RECT 83.950 18.105 84.280 18.110 ;
        RECT 89.285 18.105 89.615 18.110 ;
        RECT 94.610 18.105 94.940 18.110 ;
        RECT 99.945 18.105 100.275 18.110 ;
        RECT 105.270 18.105 105.600 18.110 ;
        RECT 110.605 18.105 110.935 18.110 ;
        RECT 115.930 18.105 116.260 18.110 ;
        RECT 121.265 18.105 121.595 18.110 ;
        RECT 126.590 18.105 126.920 18.110 ;
        RECT 29.735 16.080 30.935 16.095 ;
        RECT 31.485 16.080 31.815 16.095 ;
        RECT 36.810 16.080 37.140 16.095 ;
        RECT 42.145 16.080 42.475 16.095 ;
        RECT 47.470 16.080 47.800 16.095 ;
        RECT 52.805 16.080 53.135 16.095 ;
        RECT 58.130 16.080 58.460 16.095 ;
        RECT 63.465 16.080 63.795 16.095 ;
        RECT 68.790 16.080 69.120 16.095 ;
        RECT 74.125 16.080 74.455 16.095 ;
        RECT 79.450 16.080 79.780 16.095 ;
        RECT 84.785 16.080 85.115 16.095 ;
        RECT 90.110 16.080 90.440 16.095 ;
        RECT 95.445 16.080 95.775 16.095 ;
        RECT 100.770 16.080 101.100 16.095 ;
        RECT 106.105 16.080 106.435 16.095 ;
        RECT 111.430 16.080 111.760 16.095 ;
        RECT 116.765 16.080 117.095 16.095 ;
        RECT 122.090 16.080 122.420 16.095 ;
        RECT 29.705 15.780 127.180 16.080 ;
        RECT 29.735 15.765 30.935 15.780 ;
        RECT 31.485 15.765 31.815 15.780 ;
        RECT 36.810 15.765 37.140 15.780 ;
        RECT 42.145 15.765 42.475 15.780 ;
        RECT 47.470 15.765 47.800 15.780 ;
        RECT 52.805 15.765 53.135 15.780 ;
        RECT 58.130 15.765 58.460 15.780 ;
        RECT 63.465 15.765 63.795 15.780 ;
        RECT 68.790 15.765 69.120 15.780 ;
        RECT 74.125 15.765 74.455 15.780 ;
        RECT 79.450 15.765 79.780 15.780 ;
        RECT 84.785 15.765 85.115 15.780 ;
        RECT 90.110 15.765 90.440 15.780 ;
        RECT 95.445 15.765 95.775 15.780 ;
        RECT 100.770 15.765 101.100 15.780 ;
        RECT 106.105 15.765 106.435 15.780 ;
        RECT 111.430 15.765 111.760 15.780 ;
        RECT 116.765 15.765 117.095 15.780 ;
        RECT 122.090 15.765 122.420 15.780 ;
        RECT 29.735 15.435 30.935 15.450 ;
        RECT 35.980 15.435 36.310 15.450 ;
        RECT 41.305 15.435 41.635 15.450 ;
        RECT 46.640 15.435 46.970 15.450 ;
        RECT 51.965 15.435 52.295 15.450 ;
        RECT 57.300 15.435 57.630 15.450 ;
        RECT 62.625 15.435 62.955 15.450 ;
        RECT 67.960 15.435 68.290 15.450 ;
        RECT 73.285 15.435 73.615 15.450 ;
        RECT 78.620 15.435 78.950 15.450 ;
        RECT 83.945 15.435 84.275 15.450 ;
        RECT 89.280 15.435 89.610 15.450 ;
        RECT 94.605 15.435 94.935 15.450 ;
        RECT 99.940 15.435 100.270 15.450 ;
        RECT 105.265 15.435 105.595 15.450 ;
        RECT 110.600 15.435 110.930 15.450 ;
        RECT 115.925 15.435 116.255 15.450 ;
        RECT 121.260 15.435 121.590 15.450 ;
        RECT 126.585 15.435 126.915 15.450 ;
        RECT 29.705 15.135 127.180 15.435 ;
        RECT 29.735 15.120 30.935 15.135 ;
        RECT 35.980 15.120 36.310 15.135 ;
        RECT 41.305 15.120 41.635 15.135 ;
        RECT 46.640 15.120 46.970 15.135 ;
        RECT 51.965 15.120 52.295 15.135 ;
        RECT 57.300 15.120 57.630 15.135 ;
        RECT 62.625 15.120 62.955 15.135 ;
        RECT 67.960 15.120 68.290 15.135 ;
        RECT 73.285 15.120 73.615 15.135 ;
        RECT 78.620 15.120 78.950 15.135 ;
        RECT 83.945 15.120 84.275 15.135 ;
        RECT 89.280 15.120 89.610 15.135 ;
        RECT 94.605 15.120 94.935 15.135 ;
        RECT 99.940 15.120 100.270 15.135 ;
        RECT 105.265 15.120 105.595 15.135 ;
        RECT 110.600 15.120 110.930 15.135 ;
        RECT 115.925 15.120 116.255 15.135 ;
        RECT 121.260 15.120 121.590 15.135 ;
        RECT 126.585 15.120 126.915 15.135 ;
        RECT 29.735 14.790 30.935 14.805 ;
        RECT 31.480 14.790 31.810 14.805 ;
        RECT 36.805 14.790 37.135 14.805 ;
        RECT 42.140 14.790 42.470 14.805 ;
        RECT 47.465 14.790 47.795 14.805 ;
        RECT 52.800 14.790 53.130 14.805 ;
        RECT 58.125 14.790 58.455 14.805 ;
        RECT 63.460 14.790 63.790 14.805 ;
        RECT 68.785 14.790 69.115 14.805 ;
        RECT 74.120 14.790 74.450 14.805 ;
        RECT 79.445 14.790 79.775 14.805 ;
        RECT 84.780 14.790 85.110 14.805 ;
        RECT 90.105 14.790 90.435 14.805 ;
        RECT 95.440 14.790 95.770 14.805 ;
        RECT 100.765 14.790 101.095 14.805 ;
        RECT 106.100 14.790 106.430 14.805 ;
        RECT 111.425 14.790 111.755 14.805 ;
        RECT 116.760 14.790 117.090 14.805 ;
        RECT 122.085 14.790 122.415 14.805 ;
        RECT 29.705 14.490 127.180 14.790 ;
        RECT 29.735 14.475 30.935 14.490 ;
        RECT 31.480 14.475 31.810 14.490 ;
        RECT 36.805 14.475 37.135 14.490 ;
        RECT 42.140 14.475 42.470 14.490 ;
        RECT 47.465 14.475 47.795 14.490 ;
        RECT 52.800 14.475 53.130 14.490 ;
        RECT 58.125 14.475 58.455 14.490 ;
        RECT 63.460 14.475 63.790 14.490 ;
        RECT 68.785 14.475 69.115 14.490 ;
        RECT 74.120 14.475 74.450 14.490 ;
        RECT 79.445 14.475 79.775 14.490 ;
        RECT 84.780 14.475 85.110 14.490 ;
        RECT 90.105 14.475 90.435 14.490 ;
        RECT 95.440 14.475 95.770 14.490 ;
        RECT 100.765 14.475 101.095 14.490 ;
        RECT 106.100 14.475 106.430 14.490 ;
        RECT 111.425 14.475 111.755 14.490 ;
        RECT 116.760 14.475 117.090 14.490 ;
        RECT 122.085 14.475 122.415 14.490 ;
        RECT 29.735 14.145 30.935 14.160 ;
        RECT 35.980 14.145 36.310 14.160 ;
        RECT 41.305 14.145 41.635 14.160 ;
        RECT 46.640 14.145 46.970 14.160 ;
        RECT 51.965 14.145 52.295 14.160 ;
        RECT 57.300 14.145 57.630 14.160 ;
        RECT 62.625 14.145 62.955 14.160 ;
        RECT 67.960 14.145 68.290 14.160 ;
        RECT 73.285 14.145 73.615 14.160 ;
        RECT 78.620 14.145 78.950 14.160 ;
        RECT 83.945 14.145 84.275 14.160 ;
        RECT 89.280 14.145 89.610 14.160 ;
        RECT 94.605 14.145 94.935 14.160 ;
        RECT 99.940 14.145 100.270 14.160 ;
        RECT 105.265 14.145 105.595 14.160 ;
        RECT 110.600 14.145 110.930 14.160 ;
        RECT 115.925 14.145 116.255 14.160 ;
        RECT 121.260 14.145 121.590 14.160 ;
        RECT 126.585 14.145 126.915 14.160 ;
        RECT 29.705 13.845 127.180 14.145 ;
        RECT 29.735 13.830 30.935 13.845 ;
        RECT 35.980 13.830 36.310 13.845 ;
        RECT 41.305 13.830 41.635 13.845 ;
        RECT 46.640 13.830 46.970 13.845 ;
        RECT 51.965 13.830 52.295 13.845 ;
        RECT 57.300 13.830 57.630 13.845 ;
        RECT 62.625 13.830 62.955 13.845 ;
        RECT 67.960 13.830 68.290 13.845 ;
        RECT 73.285 13.830 73.615 13.845 ;
        RECT 78.620 13.830 78.950 13.845 ;
        RECT 83.945 13.830 84.275 13.845 ;
        RECT 89.280 13.830 89.610 13.845 ;
        RECT 94.605 13.830 94.935 13.845 ;
        RECT 99.940 13.830 100.270 13.845 ;
        RECT 105.265 13.830 105.595 13.845 ;
        RECT 110.600 13.830 110.930 13.845 ;
        RECT 115.925 13.830 116.255 13.845 ;
        RECT 121.260 13.830 121.590 13.845 ;
        RECT 126.585 13.830 126.915 13.845 ;
        RECT 29.735 12.810 30.935 12.825 ;
        RECT 31.480 12.810 31.810 12.825 ;
        RECT 36.805 12.810 37.135 12.825 ;
        RECT 42.140 12.810 42.470 12.825 ;
        RECT 47.465 12.810 47.795 12.825 ;
        RECT 52.800 12.810 53.130 12.825 ;
        RECT 58.125 12.810 58.455 12.825 ;
        RECT 63.460 12.810 63.790 12.825 ;
        RECT 68.785 12.810 69.115 12.825 ;
        RECT 74.120 12.810 74.450 12.825 ;
        RECT 79.445 12.810 79.775 12.825 ;
        RECT 84.780 12.810 85.110 12.825 ;
        RECT 90.105 12.810 90.435 12.825 ;
        RECT 95.440 12.810 95.770 12.825 ;
        RECT 100.765 12.810 101.095 12.825 ;
        RECT 106.100 12.810 106.430 12.825 ;
        RECT 111.425 12.810 111.755 12.825 ;
        RECT 116.760 12.810 117.090 12.825 ;
        RECT 122.085 12.810 122.415 12.825 ;
        RECT 29.705 12.510 127.180 12.810 ;
        RECT 29.735 12.495 30.935 12.510 ;
        RECT 31.480 12.495 31.810 12.510 ;
        RECT 36.805 12.495 37.135 12.510 ;
        RECT 42.140 12.495 42.470 12.510 ;
        RECT 47.465 12.495 47.795 12.510 ;
        RECT 52.800 12.495 53.130 12.510 ;
        RECT 58.125 12.495 58.455 12.510 ;
        RECT 63.460 12.495 63.790 12.510 ;
        RECT 68.785 12.495 69.115 12.510 ;
        RECT 74.120 12.495 74.450 12.510 ;
        RECT 79.445 12.495 79.775 12.510 ;
        RECT 84.780 12.495 85.110 12.510 ;
        RECT 90.105 12.495 90.435 12.510 ;
        RECT 95.440 12.495 95.770 12.510 ;
        RECT 100.765 12.495 101.095 12.510 ;
        RECT 106.100 12.495 106.430 12.510 ;
        RECT 111.425 12.495 111.755 12.510 ;
        RECT 116.760 12.495 117.090 12.510 ;
        RECT 122.085 12.495 122.415 12.510 ;
        RECT 29.735 12.165 30.935 12.180 ;
        RECT 35.980 12.165 36.310 12.180 ;
        RECT 41.305 12.165 41.635 12.180 ;
        RECT 46.640 12.165 46.970 12.180 ;
        RECT 51.965 12.165 52.295 12.180 ;
        RECT 57.300 12.165 57.630 12.180 ;
        RECT 62.625 12.165 62.955 12.180 ;
        RECT 67.960 12.165 68.290 12.180 ;
        RECT 73.285 12.165 73.615 12.180 ;
        RECT 78.620 12.165 78.950 12.180 ;
        RECT 83.945 12.165 84.275 12.180 ;
        RECT 89.280 12.165 89.610 12.180 ;
        RECT 94.605 12.165 94.935 12.180 ;
        RECT 99.940 12.165 100.270 12.180 ;
        RECT 105.265 12.165 105.595 12.180 ;
        RECT 110.600 12.165 110.930 12.180 ;
        RECT 115.925 12.165 116.255 12.180 ;
        RECT 121.260 12.165 121.590 12.180 ;
        RECT 126.585 12.165 126.915 12.180 ;
        RECT 29.705 11.865 127.180 12.165 ;
        RECT 29.735 11.850 30.935 11.865 ;
        RECT 35.980 11.850 36.310 11.865 ;
        RECT 41.305 11.850 41.635 11.865 ;
        RECT 46.640 11.850 46.970 11.865 ;
        RECT 51.965 11.850 52.295 11.865 ;
        RECT 57.300 11.850 57.630 11.865 ;
        RECT 62.625 11.850 62.955 11.865 ;
        RECT 67.960 11.850 68.290 11.865 ;
        RECT 73.285 11.850 73.615 11.865 ;
        RECT 78.620 11.850 78.950 11.865 ;
        RECT 83.945 11.850 84.275 11.865 ;
        RECT 89.280 11.850 89.610 11.865 ;
        RECT 94.605 11.850 94.935 11.865 ;
        RECT 99.940 11.850 100.270 11.865 ;
        RECT 105.265 11.850 105.595 11.865 ;
        RECT 110.600 11.850 110.930 11.865 ;
        RECT 115.925 11.850 116.255 11.865 ;
        RECT 121.260 11.850 121.590 11.865 ;
        RECT 126.585 11.850 126.915 11.865 ;
        RECT 29.735 11.520 30.935 11.535 ;
        RECT 31.480 11.520 31.810 11.530 ;
        RECT 36.805 11.520 37.135 11.530 ;
        RECT 42.140 11.520 42.470 11.530 ;
        RECT 47.465 11.520 47.795 11.530 ;
        RECT 52.800 11.520 53.130 11.530 ;
        RECT 58.125 11.520 58.455 11.530 ;
        RECT 63.460 11.520 63.790 11.530 ;
        RECT 68.785 11.520 69.115 11.530 ;
        RECT 74.120 11.520 74.450 11.530 ;
        RECT 79.445 11.520 79.775 11.530 ;
        RECT 84.780 11.520 85.110 11.530 ;
        RECT 90.105 11.520 90.435 11.530 ;
        RECT 95.440 11.520 95.770 11.530 ;
        RECT 100.765 11.520 101.095 11.530 ;
        RECT 106.100 11.520 106.430 11.530 ;
        RECT 111.425 11.520 111.755 11.530 ;
        RECT 116.760 11.520 117.090 11.530 ;
        RECT 122.085 11.520 122.415 11.530 ;
        RECT 29.705 11.220 127.180 11.520 ;
        RECT 29.735 11.205 30.935 11.220 ;
        RECT 31.480 11.200 31.810 11.220 ;
        RECT 36.805 11.200 37.135 11.220 ;
        RECT 42.140 11.200 42.470 11.220 ;
        RECT 47.465 11.200 47.795 11.220 ;
        RECT 52.800 11.200 53.130 11.220 ;
        RECT 58.125 11.200 58.455 11.220 ;
        RECT 63.460 11.200 63.790 11.220 ;
        RECT 68.785 11.200 69.115 11.220 ;
        RECT 74.120 11.200 74.450 11.220 ;
        RECT 79.445 11.200 79.775 11.220 ;
        RECT 84.780 11.200 85.110 11.220 ;
        RECT 90.105 11.200 90.435 11.220 ;
        RECT 95.440 11.200 95.770 11.220 ;
        RECT 100.765 11.200 101.095 11.220 ;
        RECT 106.100 11.200 106.430 11.220 ;
        RECT 111.425 11.200 111.755 11.220 ;
        RECT 116.760 11.200 117.090 11.220 ;
        RECT 122.085 11.200 122.415 11.220 ;
        RECT 29.735 10.875 30.935 10.890 ;
        RECT 35.985 10.875 36.315 10.900 ;
        RECT 41.310 10.875 41.640 10.900 ;
        RECT 46.645 10.875 46.975 10.900 ;
        RECT 51.970 10.875 52.300 10.900 ;
        RECT 57.305 10.875 57.635 10.900 ;
        RECT 62.630 10.875 62.960 10.900 ;
        RECT 67.965 10.875 68.295 10.900 ;
        RECT 73.290 10.875 73.620 10.900 ;
        RECT 78.625 10.875 78.955 10.900 ;
        RECT 83.950 10.875 84.280 10.900 ;
        RECT 89.285 10.875 89.615 10.900 ;
        RECT 94.610 10.875 94.940 10.900 ;
        RECT 99.945 10.875 100.275 10.900 ;
        RECT 105.270 10.875 105.600 10.900 ;
        RECT 110.605 10.875 110.935 10.900 ;
        RECT 115.930 10.875 116.260 10.900 ;
        RECT 121.265 10.875 121.595 10.900 ;
        RECT 126.590 10.875 126.920 10.900 ;
        RECT 29.705 10.575 127.180 10.875 ;
        RECT 29.735 10.560 30.935 10.575 ;
        RECT 35.985 10.570 36.315 10.575 ;
        RECT 41.310 10.570 41.640 10.575 ;
        RECT 46.645 10.570 46.975 10.575 ;
        RECT 51.970 10.570 52.300 10.575 ;
        RECT 57.305 10.570 57.635 10.575 ;
        RECT 62.630 10.570 62.960 10.575 ;
        RECT 67.965 10.570 68.295 10.575 ;
        RECT 73.290 10.570 73.620 10.575 ;
        RECT 78.625 10.570 78.955 10.575 ;
        RECT 83.950 10.570 84.280 10.575 ;
        RECT 89.285 10.570 89.615 10.575 ;
        RECT 94.610 10.570 94.940 10.575 ;
        RECT 99.945 10.570 100.275 10.575 ;
        RECT 105.270 10.570 105.600 10.575 ;
        RECT 110.605 10.570 110.935 10.575 ;
        RECT 115.930 10.570 116.260 10.575 ;
        RECT 121.265 10.570 121.595 10.575 ;
        RECT 126.590 10.570 126.920 10.575 ;
        RECT 38.625 9.710 39.805 10.150 ;
        RECT 44.725 9.710 45.055 9.725 ;
        RECT 38.625 9.410 45.055 9.710 ;
        RECT 38.625 8.970 39.805 9.410 ;
        RECT 44.725 9.395 45.055 9.410 ;
        RECT 49.285 9.710 50.465 10.150 ;
        RECT 55.385 9.710 55.715 9.725 ;
        RECT 49.285 9.410 55.715 9.710 ;
        RECT 49.285 8.970 50.465 9.410 ;
        RECT 55.385 9.395 55.715 9.410 ;
        RECT 59.945 9.710 61.125 10.150 ;
        RECT 66.045 9.710 66.375 9.725 ;
        RECT 59.945 9.410 66.375 9.710 ;
        RECT 59.945 8.970 61.125 9.410 ;
        RECT 66.045 9.395 66.375 9.410 ;
        RECT 70.605 9.710 71.785 10.150 ;
        RECT 76.705 9.710 77.035 9.725 ;
        RECT 70.605 9.410 77.035 9.710 ;
        RECT 70.605 8.970 71.785 9.410 ;
        RECT 76.705 9.395 77.035 9.410 ;
        RECT 81.265 9.710 82.445 10.150 ;
        RECT 87.365 9.710 87.695 9.725 ;
        RECT 81.265 9.410 87.695 9.710 ;
        RECT 81.265 8.970 82.445 9.410 ;
        RECT 87.365 9.395 87.695 9.410 ;
        RECT 91.925 9.710 93.105 10.150 ;
        RECT 98.025 9.710 98.355 9.725 ;
        RECT 91.925 9.410 98.355 9.710 ;
        RECT 91.925 8.970 93.105 9.410 ;
        RECT 98.025 9.395 98.355 9.410 ;
        RECT 102.585 9.710 103.765 10.150 ;
        RECT 108.685 9.710 109.015 9.725 ;
        RECT 102.585 9.410 109.015 9.710 ;
        RECT 102.585 8.970 103.765 9.410 ;
        RECT 108.685 9.395 109.015 9.410 ;
        RECT 113.245 9.710 114.425 10.150 ;
        RECT 119.345 9.710 119.675 9.725 ;
        RECT 113.245 9.410 119.675 9.710 ;
        RECT 113.245 8.970 114.425 9.410 ;
        RECT 119.345 9.395 119.675 9.410 ;
      LAYER met5 ;
        RECT 38.415 8.850 40.015 70.550 ;
        RECT 49.075 8.850 50.675 70.550 ;
        RECT 59.735 8.850 61.335 70.550 ;
        RECT 70.395 8.850 71.995 70.550 ;
        RECT 81.055 8.850 82.655 70.550 ;
        RECT 91.715 8.850 93.315 70.550 ;
        RECT 102.375 8.850 103.975 70.550 ;
        RECT 113.035 8.850 114.635 70.550 ;
  END
END sky130_ef_ip__rheostat_8bit
END LIBRARY

